module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
input s_162,s_163;//RE__ALLOW(00,01,10,11);
input s_164,s_165;//RE__ALLOW(00,01,10,11);
input s_166,s_167;//RE__ALLOW(00,01,10,11);
input s_168,s_169;//RE__ALLOW(00,01,10,11);
input s_170,s_171;//RE__ALLOW(00,01,10,11);
input s_172,s_173;//RE__ALLOW(00,01,10,11);
input s_174,s_175;//RE__ALLOW(00,01,10,11);
input s_176,s_177;//RE__ALLOW(00,01,10,11);
input s_178,s_179;//RE__ALLOW(00,01,10,11);
input s_180,s_181;//RE__ALLOW(00,01,10,11);
input s_182,s_183;//RE__ALLOW(00,01,10,11);
input s_184,s_185;//RE__ALLOW(00,01,10,11);
input s_186,s_187;//RE__ALLOW(00,01,10,11);
input s_188,s_189;//RE__ALLOW(00,01,10,11);
input s_190,s_191;//RE__ALLOW(00,01,10,11);
input s_192,s_193;//RE__ALLOW(00,01,10,11);
input s_194,s_195;//RE__ALLOW(00,01,10,11);
input s_196,s_197;//RE__ALLOW(00,01,10,11);
input s_198,s_199;//RE__ALLOW(00,01,10,11);
input s_200,s_201;//RE__ALLOW(00,01,10,11);
input s_202,s_203;//RE__ALLOW(00,01,10,11);
input s_204,s_205;//RE__ALLOW(00,01,10,11);
input s_206,s_207;//RE__ALLOW(00,01,10,11);
input s_208,s_209;//RE__ALLOW(00,01,10,11);
input s_210,s_211;//RE__ALLOW(00,01,10,11);
input s_212,s_213;//RE__ALLOW(00,01,10,11);
input s_214,s_215;//RE__ALLOW(00,01,10,11);
input s_216,s_217;//RE__ALLOW(00,01,10,11);
input s_218,s_219;//RE__ALLOW(00,01,10,11);
input s_220,s_221;//RE__ALLOW(00,01,10,11);
input s_222,s_223;//RE__ALLOW(00,01,10,11);
input s_224,s_225;//RE__ALLOW(00,01,10,11);
input s_226,s_227;//RE__ALLOW(00,01,10,11);
input s_228,s_229;//RE__ALLOW(00,01,10,11);
input s_230,s_231;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1499(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1500(.a(gate13inter0), .b(s_136), .O(gate13inter1));
  and2  gate1501(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1502(.a(s_136), .O(gate13inter3));
  inv1  gate1503(.a(s_137), .O(gate13inter4));
  nand2 gate1504(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1505(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1506(.a(G9), .O(gate13inter7));
  inv1  gate1507(.a(G10), .O(gate13inter8));
  nand2 gate1508(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1509(.a(s_137), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1510(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1511(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1512(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1779(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1780(.a(gate14inter0), .b(s_176), .O(gate14inter1));
  and2  gate1781(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1782(.a(s_176), .O(gate14inter3));
  inv1  gate1783(.a(s_177), .O(gate14inter4));
  nand2 gate1784(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1785(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1786(.a(G11), .O(gate14inter7));
  inv1  gate1787(.a(G12), .O(gate14inter8));
  nand2 gate1788(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1789(.a(s_177), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1790(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1791(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1792(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1625(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1626(.a(gate23inter0), .b(s_154), .O(gate23inter1));
  and2  gate1627(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1628(.a(s_154), .O(gate23inter3));
  inv1  gate1629(.a(s_155), .O(gate23inter4));
  nand2 gate1630(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1631(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1632(.a(G29), .O(gate23inter7));
  inv1  gate1633(.a(G30), .O(gate23inter8));
  nand2 gate1634(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1635(.a(s_155), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1636(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1637(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1638(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate925(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate926(.a(gate26inter0), .b(s_54), .O(gate26inter1));
  and2  gate927(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate928(.a(s_54), .O(gate26inter3));
  inv1  gate929(.a(s_55), .O(gate26inter4));
  nand2 gate930(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate931(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate932(.a(G9), .O(gate26inter7));
  inv1  gate933(.a(G13), .O(gate26inter8));
  nand2 gate934(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate935(.a(s_55), .b(gate26inter3), .O(gate26inter10));
  nor2  gate936(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate937(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate938(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1877(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1878(.a(gate31inter0), .b(s_190), .O(gate31inter1));
  and2  gate1879(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1880(.a(s_190), .O(gate31inter3));
  inv1  gate1881(.a(s_191), .O(gate31inter4));
  nand2 gate1882(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1883(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1884(.a(G4), .O(gate31inter7));
  inv1  gate1885(.a(G8), .O(gate31inter8));
  nand2 gate1886(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1887(.a(s_191), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1888(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1889(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1890(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2073(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2074(.a(gate34inter0), .b(s_218), .O(gate34inter1));
  and2  gate2075(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2076(.a(s_218), .O(gate34inter3));
  inv1  gate2077(.a(s_219), .O(gate34inter4));
  nand2 gate2078(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2079(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2080(.a(G25), .O(gate34inter7));
  inv1  gate2081(.a(G29), .O(gate34inter8));
  nand2 gate2082(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2083(.a(s_219), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2084(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2085(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2086(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate659(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate660(.a(gate43inter0), .b(s_16), .O(gate43inter1));
  and2  gate661(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate662(.a(s_16), .O(gate43inter3));
  inv1  gate663(.a(s_17), .O(gate43inter4));
  nand2 gate664(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate665(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate666(.a(G3), .O(gate43inter7));
  inv1  gate667(.a(G269), .O(gate43inter8));
  nand2 gate668(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate669(.a(s_17), .b(gate43inter3), .O(gate43inter10));
  nor2  gate670(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate671(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate672(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate799(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate800(.a(gate48inter0), .b(s_36), .O(gate48inter1));
  and2  gate801(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate802(.a(s_36), .O(gate48inter3));
  inv1  gate803(.a(s_37), .O(gate48inter4));
  nand2 gate804(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate805(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate806(.a(G8), .O(gate48inter7));
  inv1  gate807(.a(G275), .O(gate48inter8));
  nand2 gate808(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate809(.a(s_37), .b(gate48inter3), .O(gate48inter10));
  nor2  gate810(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate811(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate812(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate911(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate912(.a(gate52inter0), .b(s_52), .O(gate52inter1));
  and2  gate913(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate914(.a(s_52), .O(gate52inter3));
  inv1  gate915(.a(s_53), .O(gate52inter4));
  nand2 gate916(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate917(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate918(.a(G12), .O(gate52inter7));
  inv1  gate919(.a(G281), .O(gate52inter8));
  nand2 gate920(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate921(.a(s_53), .b(gate52inter3), .O(gate52inter10));
  nor2  gate922(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate923(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate924(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate2157(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2158(.a(gate57inter0), .b(s_230), .O(gate57inter1));
  and2  gate2159(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2160(.a(s_230), .O(gate57inter3));
  inv1  gate2161(.a(s_231), .O(gate57inter4));
  nand2 gate2162(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2163(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2164(.a(G17), .O(gate57inter7));
  inv1  gate2165(.a(G290), .O(gate57inter8));
  nand2 gate2166(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2167(.a(s_231), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2168(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2169(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2170(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2017(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2018(.a(gate59inter0), .b(s_210), .O(gate59inter1));
  and2  gate2019(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2020(.a(s_210), .O(gate59inter3));
  inv1  gate2021(.a(s_211), .O(gate59inter4));
  nand2 gate2022(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2023(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2024(.a(G19), .O(gate59inter7));
  inv1  gate2025(.a(G293), .O(gate59inter8));
  nand2 gate2026(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2027(.a(s_211), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2028(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2029(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2030(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1289(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1290(.a(gate62inter0), .b(s_106), .O(gate62inter1));
  and2  gate1291(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1292(.a(s_106), .O(gate62inter3));
  inv1  gate1293(.a(s_107), .O(gate62inter4));
  nand2 gate1294(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1295(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1296(.a(G22), .O(gate62inter7));
  inv1  gate1297(.a(G296), .O(gate62inter8));
  nand2 gate1298(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1299(.a(s_107), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1300(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1301(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1302(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1541(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1542(.a(gate64inter0), .b(s_142), .O(gate64inter1));
  and2  gate1543(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1544(.a(s_142), .O(gate64inter3));
  inv1  gate1545(.a(s_143), .O(gate64inter4));
  nand2 gate1546(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1547(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1548(.a(G24), .O(gate64inter7));
  inv1  gate1549(.a(G299), .O(gate64inter8));
  nand2 gate1550(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1551(.a(s_143), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1552(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1553(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1554(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate2045(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2046(.a(gate65inter0), .b(s_214), .O(gate65inter1));
  and2  gate2047(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2048(.a(s_214), .O(gate65inter3));
  inv1  gate2049(.a(s_215), .O(gate65inter4));
  nand2 gate2050(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2051(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2052(.a(G25), .O(gate65inter7));
  inv1  gate2053(.a(G302), .O(gate65inter8));
  nand2 gate2054(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2055(.a(s_215), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2056(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2057(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2058(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1989(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1990(.a(gate66inter0), .b(s_206), .O(gate66inter1));
  and2  gate1991(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1992(.a(s_206), .O(gate66inter3));
  inv1  gate1993(.a(s_207), .O(gate66inter4));
  nand2 gate1994(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1995(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1996(.a(G26), .O(gate66inter7));
  inv1  gate1997(.a(G302), .O(gate66inter8));
  nand2 gate1998(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1999(.a(s_207), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2000(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2001(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2002(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1709(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1710(.a(gate70inter0), .b(s_166), .O(gate70inter1));
  and2  gate1711(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1712(.a(s_166), .O(gate70inter3));
  inv1  gate1713(.a(s_167), .O(gate70inter4));
  nand2 gate1714(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1715(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1716(.a(G30), .O(gate70inter7));
  inv1  gate1717(.a(G308), .O(gate70inter8));
  nand2 gate1718(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1719(.a(s_167), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1720(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1721(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1722(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1849(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1850(.a(gate72inter0), .b(s_186), .O(gate72inter1));
  and2  gate1851(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1852(.a(s_186), .O(gate72inter3));
  inv1  gate1853(.a(s_187), .O(gate72inter4));
  nand2 gate1854(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1855(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1856(.a(G32), .O(gate72inter7));
  inv1  gate1857(.a(G311), .O(gate72inter8));
  nand2 gate1858(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1859(.a(s_187), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1860(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1861(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1862(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1443(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1444(.a(gate73inter0), .b(s_128), .O(gate73inter1));
  and2  gate1445(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1446(.a(s_128), .O(gate73inter3));
  inv1  gate1447(.a(s_129), .O(gate73inter4));
  nand2 gate1448(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1449(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1450(.a(G1), .O(gate73inter7));
  inv1  gate1451(.a(G314), .O(gate73inter8));
  nand2 gate1452(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1453(.a(s_129), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1454(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1455(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1456(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate2101(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2102(.a(gate81inter0), .b(s_222), .O(gate81inter1));
  and2  gate2103(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2104(.a(s_222), .O(gate81inter3));
  inv1  gate2105(.a(s_223), .O(gate81inter4));
  nand2 gate2106(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2107(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2108(.a(G3), .O(gate81inter7));
  inv1  gate2109(.a(G326), .O(gate81inter8));
  nand2 gate2110(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2111(.a(s_223), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2112(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2113(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2114(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1527(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1528(.a(gate82inter0), .b(s_140), .O(gate82inter1));
  and2  gate1529(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1530(.a(s_140), .O(gate82inter3));
  inv1  gate1531(.a(s_141), .O(gate82inter4));
  nand2 gate1532(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1533(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1534(.a(G7), .O(gate82inter7));
  inv1  gate1535(.a(G326), .O(gate82inter8));
  nand2 gate1536(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1537(.a(s_141), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1538(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1539(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1540(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1429(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1430(.a(gate85inter0), .b(s_126), .O(gate85inter1));
  and2  gate1431(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1432(.a(s_126), .O(gate85inter3));
  inv1  gate1433(.a(s_127), .O(gate85inter4));
  nand2 gate1434(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1435(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1436(.a(G4), .O(gate85inter7));
  inv1  gate1437(.a(G332), .O(gate85inter8));
  nand2 gate1438(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1439(.a(s_127), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1440(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1441(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1442(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1415(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1416(.a(gate86inter0), .b(s_124), .O(gate86inter1));
  and2  gate1417(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1418(.a(s_124), .O(gate86inter3));
  inv1  gate1419(.a(s_125), .O(gate86inter4));
  nand2 gate1420(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1421(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1422(.a(G8), .O(gate86inter7));
  inv1  gate1423(.a(G332), .O(gate86inter8));
  nand2 gate1424(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1425(.a(s_125), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1426(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1427(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1428(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate589(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate590(.a(gate88inter0), .b(s_6), .O(gate88inter1));
  and2  gate591(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate592(.a(s_6), .O(gate88inter3));
  inv1  gate593(.a(s_7), .O(gate88inter4));
  nand2 gate594(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate595(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate596(.a(G16), .O(gate88inter7));
  inv1  gate597(.a(G335), .O(gate88inter8));
  nand2 gate598(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate599(.a(s_7), .b(gate88inter3), .O(gate88inter10));
  nor2  gate600(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate601(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate602(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate1471(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1472(.a(gate89inter0), .b(s_132), .O(gate89inter1));
  and2  gate1473(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1474(.a(s_132), .O(gate89inter3));
  inv1  gate1475(.a(s_133), .O(gate89inter4));
  nand2 gate1476(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1477(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1478(.a(G17), .O(gate89inter7));
  inv1  gate1479(.a(G338), .O(gate89inter8));
  nand2 gate1480(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1481(.a(s_133), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1482(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1483(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1484(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1317(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1318(.a(gate92inter0), .b(s_110), .O(gate92inter1));
  and2  gate1319(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1320(.a(s_110), .O(gate92inter3));
  inv1  gate1321(.a(s_111), .O(gate92inter4));
  nand2 gate1322(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1323(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1324(.a(G29), .O(gate92inter7));
  inv1  gate1325(.a(G341), .O(gate92inter8));
  nand2 gate1326(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1327(.a(s_111), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1328(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1329(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1330(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate575(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate576(.a(gate94inter0), .b(s_4), .O(gate94inter1));
  and2  gate577(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate578(.a(s_4), .O(gate94inter3));
  inv1  gate579(.a(s_5), .O(gate94inter4));
  nand2 gate580(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate581(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate582(.a(G22), .O(gate94inter7));
  inv1  gate583(.a(G344), .O(gate94inter8));
  nand2 gate584(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate585(.a(s_5), .b(gate94inter3), .O(gate94inter10));
  nor2  gate586(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate587(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate588(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate1485(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1486(.a(gate95inter0), .b(s_134), .O(gate95inter1));
  and2  gate1487(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1488(.a(s_134), .O(gate95inter3));
  inv1  gate1489(.a(s_135), .O(gate95inter4));
  nand2 gate1490(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1491(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1492(.a(G26), .O(gate95inter7));
  inv1  gate1493(.a(G347), .O(gate95inter8));
  nand2 gate1494(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1495(.a(s_135), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1496(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1497(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1498(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate939(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate940(.a(gate98inter0), .b(s_56), .O(gate98inter1));
  and2  gate941(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate942(.a(s_56), .O(gate98inter3));
  inv1  gate943(.a(s_57), .O(gate98inter4));
  nand2 gate944(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate945(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate946(.a(G23), .O(gate98inter7));
  inv1  gate947(.a(G350), .O(gate98inter8));
  nand2 gate948(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate949(.a(s_57), .b(gate98inter3), .O(gate98inter10));
  nor2  gate950(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate951(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate952(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1751(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1752(.a(gate105inter0), .b(s_172), .O(gate105inter1));
  and2  gate1753(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1754(.a(s_172), .O(gate105inter3));
  inv1  gate1755(.a(s_173), .O(gate105inter4));
  nand2 gate1756(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1757(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1758(.a(G362), .O(gate105inter7));
  inv1  gate1759(.a(G363), .O(gate105inter8));
  nand2 gate1760(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1761(.a(s_173), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1762(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1763(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1764(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1639(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1640(.a(gate107inter0), .b(s_156), .O(gate107inter1));
  and2  gate1641(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1642(.a(s_156), .O(gate107inter3));
  inv1  gate1643(.a(s_157), .O(gate107inter4));
  nand2 gate1644(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1645(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1646(.a(G366), .O(gate107inter7));
  inv1  gate1647(.a(G367), .O(gate107inter8));
  nand2 gate1648(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1649(.a(s_157), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1650(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1651(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1652(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1919(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1920(.a(gate114inter0), .b(s_196), .O(gate114inter1));
  and2  gate1921(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1922(.a(s_196), .O(gate114inter3));
  inv1  gate1923(.a(s_197), .O(gate114inter4));
  nand2 gate1924(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1925(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1926(.a(G380), .O(gate114inter7));
  inv1  gate1927(.a(G381), .O(gate114inter8));
  nand2 gate1928(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1929(.a(s_197), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1930(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1931(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1932(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1079(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1080(.a(gate116inter0), .b(s_76), .O(gate116inter1));
  and2  gate1081(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1082(.a(s_76), .O(gate116inter3));
  inv1  gate1083(.a(s_77), .O(gate116inter4));
  nand2 gate1084(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1085(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1086(.a(G384), .O(gate116inter7));
  inv1  gate1087(.a(G385), .O(gate116inter8));
  nand2 gate1088(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1089(.a(s_77), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1090(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1091(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1092(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1023(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1024(.a(gate124inter0), .b(s_68), .O(gate124inter1));
  and2  gate1025(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1026(.a(s_68), .O(gate124inter3));
  inv1  gate1027(.a(s_69), .O(gate124inter4));
  nand2 gate1028(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1029(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1030(.a(G400), .O(gate124inter7));
  inv1  gate1031(.a(G401), .O(gate124inter8));
  nand2 gate1032(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1033(.a(s_69), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1034(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1035(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1036(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate2087(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2088(.a(gate125inter0), .b(s_220), .O(gate125inter1));
  and2  gate2089(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2090(.a(s_220), .O(gate125inter3));
  inv1  gate2091(.a(s_221), .O(gate125inter4));
  nand2 gate2092(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2093(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2094(.a(G402), .O(gate125inter7));
  inv1  gate2095(.a(G403), .O(gate125inter8));
  nand2 gate2096(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2097(.a(s_221), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2098(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2099(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2100(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate1009(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1010(.a(gate131inter0), .b(s_66), .O(gate131inter1));
  and2  gate1011(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1012(.a(s_66), .O(gate131inter3));
  inv1  gate1013(.a(s_67), .O(gate131inter4));
  nand2 gate1014(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1015(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1016(.a(G414), .O(gate131inter7));
  inv1  gate1017(.a(G415), .O(gate131inter8));
  nand2 gate1018(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1019(.a(s_67), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1020(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1021(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1022(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate687(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate688(.a(gate137inter0), .b(s_20), .O(gate137inter1));
  and2  gate689(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate690(.a(s_20), .O(gate137inter3));
  inv1  gate691(.a(s_21), .O(gate137inter4));
  nand2 gate692(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate693(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate694(.a(G426), .O(gate137inter7));
  inv1  gate695(.a(G429), .O(gate137inter8));
  nand2 gate696(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate697(.a(s_21), .b(gate137inter3), .O(gate137inter10));
  nor2  gate698(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate699(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate700(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1555(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1556(.a(gate139inter0), .b(s_144), .O(gate139inter1));
  and2  gate1557(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1558(.a(s_144), .O(gate139inter3));
  inv1  gate1559(.a(s_145), .O(gate139inter4));
  nand2 gate1560(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1561(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1562(.a(G438), .O(gate139inter7));
  inv1  gate1563(.a(G441), .O(gate139inter8));
  nand2 gate1564(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1565(.a(s_145), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1566(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1567(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1568(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1765(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1766(.a(gate140inter0), .b(s_174), .O(gate140inter1));
  and2  gate1767(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1768(.a(s_174), .O(gate140inter3));
  inv1  gate1769(.a(s_175), .O(gate140inter4));
  nand2 gate1770(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1771(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1772(.a(G444), .O(gate140inter7));
  inv1  gate1773(.a(G447), .O(gate140inter8));
  nand2 gate1774(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1775(.a(s_175), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1776(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1777(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1778(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1835(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1836(.a(gate142inter0), .b(s_184), .O(gate142inter1));
  and2  gate1837(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1838(.a(s_184), .O(gate142inter3));
  inv1  gate1839(.a(s_185), .O(gate142inter4));
  nand2 gate1840(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1841(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1842(.a(G456), .O(gate142inter7));
  inv1  gate1843(.a(G459), .O(gate142inter8));
  nand2 gate1844(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1845(.a(s_185), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1846(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1847(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1848(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1401(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1402(.a(gate144inter0), .b(s_122), .O(gate144inter1));
  and2  gate1403(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1404(.a(s_122), .O(gate144inter3));
  inv1  gate1405(.a(s_123), .O(gate144inter4));
  nand2 gate1406(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1407(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1408(.a(G468), .O(gate144inter7));
  inv1  gate1409(.a(G471), .O(gate144inter8));
  nand2 gate1410(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1411(.a(s_123), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1412(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1413(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1414(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate729(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate730(.a(gate147inter0), .b(s_26), .O(gate147inter1));
  and2  gate731(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate732(.a(s_26), .O(gate147inter3));
  inv1  gate733(.a(s_27), .O(gate147inter4));
  nand2 gate734(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate735(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate736(.a(G486), .O(gate147inter7));
  inv1  gate737(.a(G489), .O(gate147inter8));
  nand2 gate738(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate739(.a(s_27), .b(gate147inter3), .O(gate147inter10));
  nor2  gate740(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate741(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate742(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1891(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1892(.a(gate150inter0), .b(s_192), .O(gate150inter1));
  and2  gate1893(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1894(.a(s_192), .O(gate150inter3));
  inv1  gate1895(.a(s_193), .O(gate150inter4));
  nand2 gate1896(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1897(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1898(.a(G504), .O(gate150inter7));
  inv1  gate1899(.a(G507), .O(gate150inter8));
  nand2 gate1900(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1901(.a(s_193), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1902(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1903(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1904(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate995(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate996(.a(gate155inter0), .b(s_64), .O(gate155inter1));
  and2  gate997(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate998(.a(s_64), .O(gate155inter3));
  inv1  gate999(.a(s_65), .O(gate155inter4));
  nand2 gate1000(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1001(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1002(.a(G432), .O(gate155inter7));
  inv1  gate1003(.a(G525), .O(gate155inter8));
  nand2 gate1004(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1005(.a(s_65), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1006(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1007(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1008(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate841(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate842(.a(gate159inter0), .b(s_42), .O(gate159inter1));
  and2  gate843(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate844(.a(s_42), .O(gate159inter3));
  inv1  gate845(.a(s_43), .O(gate159inter4));
  nand2 gate846(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate847(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate848(.a(G444), .O(gate159inter7));
  inv1  gate849(.a(G531), .O(gate159inter8));
  nand2 gate850(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate851(.a(s_43), .b(gate159inter3), .O(gate159inter10));
  nor2  gate852(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate853(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate854(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1653(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1654(.a(gate168inter0), .b(s_158), .O(gate168inter1));
  and2  gate1655(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1656(.a(s_158), .O(gate168inter3));
  inv1  gate1657(.a(s_159), .O(gate168inter4));
  nand2 gate1658(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1659(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1660(.a(G471), .O(gate168inter7));
  inv1  gate1661(.a(G543), .O(gate168inter8));
  nand2 gate1662(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1663(.a(s_159), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1664(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1665(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1666(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1191(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1192(.a(gate169inter0), .b(s_92), .O(gate169inter1));
  and2  gate1193(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1194(.a(s_92), .O(gate169inter3));
  inv1  gate1195(.a(s_93), .O(gate169inter4));
  nand2 gate1196(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1197(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1198(.a(G474), .O(gate169inter7));
  inv1  gate1199(.a(G546), .O(gate169inter8));
  nand2 gate1200(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1201(.a(s_93), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1202(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1203(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1204(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1359(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1360(.a(gate170inter0), .b(s_116), .O(gate170inter1));
  and2  gate1361(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1362(.a(s_116), .O(gate170inter3));
  inv1  gate1363(.a(s_117), .O(gate170inter4));
  nand2 gate1364(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1365(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1366(.a(G477), .O(gate170inter7));
  inv1  gate1367(.a(G546), .O(gate170inter8));
  nand2 gate1368(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1369(.a(s_117), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1370(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1371(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1372(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1569(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1570(.a(gate174inter0), .b(s_146), .O(gate174inter1));
  and2  gate1571(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1572(.a(s_146), .O(gate174inter3));
  inv1  gate1573(.a(s_147), .O(gate174inter4));
  nand2 gate1574(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1575(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1576(.a(G489), .O(gate174inter7));
  inv1  gate1577(.a(G552), .O(gate174inter8));
  nand2 gate1578(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1579(.a(s_147), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1580(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1581(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1582(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1793(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1794(.a(gate175inter0), .b(s_178), .O(gate175inter1));
  and2  gate1795(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1796(.a(s_178), .O(gate175inter3));
  inv1  gate1797(.a(s_179), .O(gate175inter4));
  nand2 gate1798(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1799(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1800(.a(G492), .O(gate175inter7));
  inv1  gate1801(.a(G555), .O(gate175inter8));
  nand2 gate1802(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1803(.a(s_179), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1804(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1805(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1806(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate561(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate562(.a(gate179inter0), .b(s_2), .O(gate179inter1));
  and2  gate563(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate564(.a(s_2), .O(gate179inter3));
  inv1  gate565(.a(s_3), .O(gate179inter4));
  nand2 gate566(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate567(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate568(.a(G504), .O(gate179inter7));
  inv1  gate569(.a(G561), .O(gate179inter8));
  nand2 gate570(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate571(.a(s_3), .b(gate179inter3), .O(gate179inter10));
  nor2  gate572(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate573(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate574(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1611(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1612(.a(gate180inter0), .b(s_152), .O(gate180inter1));
  and2  gate1613(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1614(.a(s_152), .O(gate180inter3));
  inv1  gate1615(.a(s_153), .O(gate180inter4));
  nand2 gate1616(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1617(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1618(.a(G507), .O(gate180inter7));
  inv1  gate1619(.a(G561), .O(gate180inter8));
  nand2 gate1620(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1621(.a(s_153), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1622(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1623(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1624(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1135(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1136(.a(gate186inter0), .b(s_84), .O(gate186inter1));
  and2  gate1137(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1138(.a(s_84), .O(gate186inter3));
  inv1  gate1139(.a(s_85), .O(gate186inter4));
  nand2 gate1140(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1141(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1142(.a(G572), .O(gate186inter7));
  inv1  gate1143(.a(G573), .O(gate186inter8));
  nand2 gate1144(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1145(.a(s_85), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1146(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1147(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1148(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate631(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate632(.a(gate187inter0), .b(s_12), .O(gate187inter1));
  and2  gate633(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate634(.a(s_12), .O(gate187inter3));
  inv1  gate635(.a(s_13), .O(gate187inter4));
  nand2 gate636(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate637(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate638(.a(G574), .O(gate187inter7));
  inv1  gate639(.a(G575), .O(gate187inter8));
  nand2 gate640(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate641(.a(s_13), .b(gate187inter3), .O(gate187inter10));
  nor2  gate642(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate643(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate644(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1961(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1962(.a(gate188inter0), .b(s_202), .O(gate188inter1));
  and2  gate1963(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1964(.a(s_202), .O(gate188inter3));
  inv1  gate1965(.a(s_203), .O(gate188inter4));
  nand2 gate1966(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1967(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1968(.a(G576), .O(gate188inter7));
  inv1  gate1969(.a(G577), .O(gate188inter8));
  nand2 gate1970(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1971(.a(s_203), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1972(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1973(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1974(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1233(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1234(.a(gate190inter0), .b(s_98), .O(gate190inter1));
  and2  gate1235(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1236(.a(s_98), .O(gate190inter3));
  inv1  gate1237(.a(s_99), .O(gate190inter4));
  nand2 gate1238(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1239(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1240(.a(G580), .O(gate190inter7));
  inv1  gate1241(.a(G581), .O(gate190inter8));
  nand2 gate1242(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1243(.a(s_99), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1244(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1245(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1246(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2003(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2004(.a(gate191inter0), .b(s_208), .O(gate191inter1));
  and2  gate2005(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2006(.a(s_208), .O(gate191inter3));
  inv1  gate2007(.a(s_209), .O(gate191inter4));
  nand2 gate2008(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2009(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2010(.a(G582), .O(gate191inter7));
  inv1  gate2011(.a(G583), .O(gate191inter8));
  nand2 gate2012(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2013(.a(s_209), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2014(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2015(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2016(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1723(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1724(.a(gate192inter0), .b(s_168), .O(gate192inter1));
  and2  gate1725(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1726(.a(s_168), .O(gate192inter3));
  inv1  gate1727(.a(s_169), .O(gate192inter4));
  nand2 gate1728(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1729(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1730(.a(G584), .O(gate192inter7));
  inv1  gate1731(.a(G585), .O(gate192inter8));
  nand2 gate1732(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1733(.a(s_169), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1734(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1735(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1736(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1247(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1248(.a(gate195inter0), .b(s_100), .O(gate195inter1));
  and2  gate1249(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1250(.a(s_100), .O(gate195inter3));
  inv1  gate1251(.a(s_101), .O(gate195inter4));
  nand2 gate1252(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1253(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1254(.a(G590), .O(gate195inter7));
  inv1  gate1255(.a(G591), .O(gate195inter8));
  nand2 gate1256(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1257(.a(s_101), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1258(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1259(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1260(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2129(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2130(.a(gate200inter0), .b(s_226), .O(gate200inter1));
  and2  gate2131(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2132(.a(s_226), .O(gate200inter3));
  inv1  gate2133(.a(s_227), .O(gate200inter4));
  nand2 gate2134(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2135(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2136(.a(G600), .O(gate200inter7));
  inv1  gate2137(.a(G601), .O(gate200inter8));
  nand2 gate2138(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2139(.a(s_227), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2140(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2141(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2142(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1219(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1220(.a(gate229inter0), .b(s_96), .O(gate229inter1));
  and2  gate1221(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1222(.a(s_96), .O(gate229inter3));
  inv1  gate1223(.a(s_97), .O(gate229inter4));
  nand2 gate1224(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1225(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1226(.a(G698), .O(gate229inter7));
  inv1  gate1227(.a(G699), .O(gate229inter8));
  nand2 gate1228(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1229(.a(s_97), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1230(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1231(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1232(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1947(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1948(.a(gate231inter0), .b(s_200), .O(gate231inter1));
  and2  gate1949(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1950(.a(s_200), .O(gate231inter3));
  inv1  gate1951(.a(s_201), .O(gate231inter4));
  nand2 gate1952(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1953(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1954(.a(G702), .O(gate231inter7));
  inv1  gate1955(.a(G703), .O(gate231inter8));
  nand2 gate1956(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1957(.a(s_201), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1958(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1959(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1960(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1037(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1038(.a(gate232inter0), .b(s_70), .O(gate232inter1));
  and2  gate1039(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1040(.a(s_70), .O(gate232inter3));
  inv1  gate1041(.a(s_71), .O(gate232inter4));
  nand2 gate1042(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1043(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1044(.a(G704), .O(gate232inter7));
  inv1  gate1045(.a(G705), .O(gate232inter8));
  nand2 gate1046(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1047(.a(s_71), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1048(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1049(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1050(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1163(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1164(.a(gate238inter0), .b(s_88), .O(gate238inter1));
  and2  gate1165(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1166(.a(s_88), .O(gate238inter3));
  inv1  gate1167(.a(s_89), .O(gate238inter4));
  nand2 gate1168(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1169(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1170(.a(G257), .O(gate238inter7));
  inv1  gate1171(.a(G709), .O(gate238inter8));
  nand2 gate1172(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1173(.a(s_89), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1174(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1175(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1176(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1821(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1822(.a(gate241inter0), .b(s_182), .O(gate241inter1));
  and2  gate1823(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1824(.a(s_182), .O(gate241inter3));
  inv1  gate1825(.a(s_183), .O(gate241inter4));
  nand2 gate1826(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1827(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1828(.a(G242), .O(gate241inter7));
  inv1  gate1829(.a(G730), .O(gate241inter8));
  nand2 gate1830(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1831(.a(s_183), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1832(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1833(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1834(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1695(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1696(.a(gate245inter0), .b(s_164), .O(gate245inter1));
  and2  gate1697(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1698(.a(s_164), .O(gate245inter3));
  inv1  gate1699(.a(s_165), .O(gate245inter4));
  nand2 gate1700(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1701(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1702(.a(G248), .O(gate245inter7));
  inv1  gate1703(.a(G736), .O(gate245inter8));
  nand2 gate1704(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1705(.a(s_165), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1706(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1707(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1708(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate1149(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1150(.a(gate246inter0), .b(s_86), .O(gate246inter1));
  and2  gate1151(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1152(.a(s_86), .O(gate246inter3));
  inv1  gate1153(.a(s_87), .O(gate246inter4));
  nand2 gate1154(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1155(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1156(.a(G724), .O(gate246inter7));
  inv1  gate1157(.a(G736), .O(gate246inter8));
  nand2 gate1158(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1159(.a(s_87), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1160(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1161(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1162(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate897(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate898(.a(gate248inter0), .b(s_50), .O(gate248inter1));
  and2  gate899(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate900(.a(s_50), .O(gate248inter3));
  inv1  gate901(.a(s_51), .O(gate248inter4));
  nand2 gate902(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate903(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate904(.a(G727), .O(gate248inter7));
  inv1  gate905(.a(G739), .O(gate248inter8));
  nand2 gate906(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate907(.a(s_51), .b(gate248inter3), .O(gate248inter10));
  nor2  gate908(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate909(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate910(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate701(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate702(.a(gate253inter0), .b(s_22), .O(gate253inter1));
  and2  gate703(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate704(.a(s_22), .O(gate253inter3));
  inv1  gate705(.a(s_23), .O(gate253inter4));
  nand2 gate706(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate707(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate708(.a(G260), .O(gate253inter7));
  inv1  gate709(.a(G748), .O(gate253inter8));
  nand2 gate710(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate711(.a(s_23), .b(gate253inter3), .O(gate253inter10));
  nor2  gate712(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate713(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate714(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1513(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1514(.a(gate260inter0), .b(s_138), .O(gate260inter1));
  and2  gate1515(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1516(.a(s_138), .O(gate260inter3));
  inv1  gate1517(.a(s_139), .O(gate260inter4));
  nand2 gate1518(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1519(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1520(.a(G760), .O(gate260inter7));
  inv1  gate1521(.a(G761), .O(gate260inter8));
  nand2 gate1522(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1523(.a(s_139), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1524(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1525(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1526(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1933(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1934(.a(gate262inter0), .b(s_198), .O(gate262inter1));
  and2  gate1935(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1936(.a(s_198), .O(gate262inter3));
  inv1  gate1937(.a(s_199), .O(gate262inter4));
  nand2 gate1938(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1939(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1940(.a(G764), .O(gate262inter7));
  inv1  gate1941(.a(G765), .O(gate262inter8));
  nand2 gate1942(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1943(.a(s_199), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1944(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1945(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1946(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1107(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1108(.a(gate274inter0), .b(s_80), .O(gate274inter1));
  and2  gate1109(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1110(.a(s_80), .O(gate274inter3));
  inv1  gate1111(.a(s_81), .O(gate274inter4));
  nand2 gate1112(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1113(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1114(.a(G770), .O(gate274inter7));
  inv1  gate1115(.a(G794), .O(gate274inter8));
  nand2 gate1116(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1117(.a(s_81), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1118(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1119(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1120(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate953(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate954(.a(gate277inter0), .b(s_58), .O(gate277inter1));
  and2  gate955(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate956(.a(s_58), .O(gate277inter3));
  inv1  gate957(.a(s_59), .O(gate277inter4));
  nand2 gate958(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate959(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate960(.a(G648), .O(gate277inter7));
  inv1  gate961(.a(G800), .O(gate277inter8));
  nand2 gate962(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate963(.a(s_59), .b(gate277inter3), .O(gate277inter10));
  nor2  gate964(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate965(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate966(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate869(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate870(.a(gate281inter0), .b(s_46), .O(gate281inter1));
  and2  gate871(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate872(.a(s_46), .O(gate281inter3));
  inv1  gate873(.a(s_47), .O(gate281inter4));
  nand2 gate874(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate875(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate876(.a(G654), .O(gate281inter7));
  inv1  gate877(.a(G806), .O(gate281inter8));
  nand2 gate878(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate879(.a(s_47), .b(gate281inter3), .O(gate281inter10));
  nor2  gate880(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate881(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate882(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1205(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1206(.a(gate290inter0), .b(s_94), .O(gate290inter1));
  and2  gate1207(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1208(.a(s_94), .O(gate290inter3));
  inv1  gate1209(.a(s_95), .O(gate290inter4));
  nand2 gate1210(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1211(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1212(.a(G820), .O(gate290inter7));
  inv1  gate1213(.a(G821), .O(gate290inter8));
  nand2 gate1214(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1215(.a(s_95), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1216(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1217(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1218(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate547(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate548(.a(gate293inter0), .b(s_0), .O(gate293inter1));
  and2  gate549(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate550(.a(s_0), .O(gate293inter3));
  inv1  gate551(.a(s_1), .O(gate293inter4));
  nand2 gate552(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate553(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate554(.a(G828), .O(gate293inter7));
  inv1  gate555(.a(G829), .O(gate293inter8));
  nand2 gate556(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate557(.a(s_1), .b(gate293inter3), .O(gate293inter10));
  nor2  gate558(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate559(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate560(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1065(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1066(.a(gate294inter0), .b(s_74), .O(gate294inter1));
  and2  gate1067(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1068(.a(s_74), .O(gate294inter3));
  inv1  gate1069(.a(s_75), .O(gate294inter4));
  nand2 gate1070(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1071(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1072(.a(G832), .O(gate294inter7));
  inv1  gate1073(.a(G833), .O(gate294inter8));
  nand2 gate1074(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1075(.a(s_75), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1076(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1077(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1078(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1387(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1388(.a(gate296inter0), .b(s_120), .O(gate296inter1));
  and2  gate1389(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1390(.a(s_120), .O(gate296inter3));
  inv1  gate1391(.a(s_121), .O(gate296inter4));
  nand2 gate1392(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1393(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1394(.a(G826), .O(gate296inter7));
  inv1  gate1395(.a(G827), .O(gate296inter8));
  nand2 gate1396(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1397(.a(s_121), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1398(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1399(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1400(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1303(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1304(.a(gate388inter0), .b(s_108), .O(gate388inter1));
  and2  gate1305(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1306(.a(s_108), .O(gate388inter3));
  inv1  gate1307(.a(s_109), .O(gate388inter4));
  nand2 gate1308(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1309(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1310(.a(G2), .O(gate388inter7));
  inv1  gate1311(.a(G1039), .O(gate388inter8));
  nand2 gate1312(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1313(.a(s_109), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1314(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1315(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1316(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1051(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1052(.a(gate393inter0), .b(s_72), .O(gate393inter1));
  and2  gate1053(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1054(.a(s_72), .O(gate393inter3));
  inv1  gate1055(.a(s_73), .O(gate393inter4));
  nand2 gate1056(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1057(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1058(.a(G7), .O(gate393inter7));
  inv1  gate1059(.a(G1054), .O(gate393inter8));
  nand2 gate1060(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1061(.a(s_73), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1062(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1063(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1064(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1905(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1906(.a(gate398inter0), .b(s_194), .O(gate398inter1));
  and2  gate1907(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1908(.a(s_194), .O(gate398inter3));
  inv1  gate1909(.a(s_195), .O(gate398inter4));
  nand2 gate1910(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1911(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1912(.a(G12), .O(gate398inter7));
  inv1  gate1913(.a(G1069), .O(gate398inter8));
  nand2 gate1914(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1915(.a(s_195), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1916(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1917(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1918(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1457(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1458(.a(gate406inter0), .b(s_130), .O(gate406inter1));
  and2  gate1459(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1460(.a(s_130), .O(gate406inter3));
  inv1  gate1461(.a(s_131), .O(gate406inter4));
  nand2 gate1462(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1463(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1464(.a(G20), .O(gate406inter7));
  inv1  gate1465(.a(G1093), .O(gate406inter8));
  nand2 gate1466(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1467(.a(s_131), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1468(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1469(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1470(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate981(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate982(.a(gate407inter0), .b(s_62), .O(gate407inter1));
  and2  gate983(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate984(.a(s_62), .O(gate407inter3));
  inv1  gate985(.a(s_63), .O(gate407inter4));
  nand2 gate986(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate987(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate988(.a(G21), .O(gate407inter7));
  inv1  gate989(.a(G1096), .O(gate407inter8));
  nand2 gate990(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate991(.a(s_63), .b(gate407inter3), .O(gate407inter10));
  nor2  gate992(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate993(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate994(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1373(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1374(.a(gate409inter0), .b(s_118), .O(gate409inter1));
  and2  gate1375(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1376(.a(s_118), .O(gate409inter3));
  inv1  gate1377(.a(s_119), .O(gate409inter4));
  nand2 gate1378(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1379(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1380(.a(G23), .O(gate409inter7));
  inv1  gate1381(.a(G1102), .O(gate409inter8));
  nand2 gate1382(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1383(.a(s_119), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1384(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1385(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1386(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2115(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2116(.a(gate411inter0), .b(s_224), .O(gate411inter1));
  and2  gate2117(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2118(.a(s_224), .O(gate411inter3));
  inv1  gate2119(.a(s_225), .O(gate411inter4));
  nand2 gate2120(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2121(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2122(.a(G25), .O(gate411inter7));
  inv1  gate2123(.a(G1108), .O(gate411inter8));
  nand2 gate2124(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2125(.a(s_225), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2126(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2127(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2128(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1093(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1094(.a(gate415inter0), .b(s_78), .O(gate415inter1));
  and2  gate1095(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1096(.a(s_78), .O(gate415inter3));
  inv1  gate1097(.a(s_79), .O(gate415inter4));
  nand2 gate1098(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1099(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1100(.a(G29), .O(gate415inter7));
  inv1  gate1101(.a(G1120), .O(gate415inter8));
  nand2 gate1102(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1103(.a(s_79), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1104(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1105(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1106(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1737(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1738(.a(gate420inter0), .b(s_170), .O(gate420inter1));
  and2  gate1739(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1740(.a(s_170), .O(gate420inter3));
  inv1  gate1741(.a(s_171), .O(gate420inter4));
  nand2 gate1742(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1743(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1744(.a(G1036), .O(gate420inter7));
  inv1  gate1745(.a(G1132), .O(gate420inter8));
  nand2 gate1746(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1747(.a(s_171), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1748(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1749(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1750(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1807(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1808(.a(gate423inter0), .b(s_180), .O(gate423inter1));
  and2  gate1809(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1810(.a(s_180), .O(gate423inter3));
  inv1  gate1811(.a(s_181), .O(gate423inter4));
  nand2 gate1812(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1813(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1814(.a(G3), .O(gate423inter7));
  inv1  gate1815(.a(G1138), .O(gate423inter8));
  nand2 gate1816(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1817(.a(s_181), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1818(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1819(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1820(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1261(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1262(.a(gate426inter0), .b(s_102), .O(gate426inter1));
  and2  gate1263(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1264(.a(s_102), .O(gate426inter3));
  inv1  gate1265(.a(s_103), .O(gate426inter4));
  nand2 gate1266(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1267(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1268(.a(G1045), .O(gate426inter7));
  inv1  gate1269(.a(G1141), .O(gate426inter8));
  nand2 gate1270(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1271(.a(s_103), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1272(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1273(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1274(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2059(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2060(.a(gate427inter0), .b(s_216), .O(gate427inter1));
  and2  gate2061(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2062(.a(s_216), .O(gate427inter3));
  inv1  gate2063(.a(s_217), .O(gate427inter4));
  nand2 gate2064(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2065(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2066(.a(G5), .O(gate427inter7));
  inv1  gate2067(.a(G1144), .O(gate427inter8));
  nand2 gate2068(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2069(.a(s_217), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2070(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2071(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2072(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate967(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate968(.a(gate428inter0), .b(s_60), .O(gate428inter1));
  and2  gate969(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate970(.a(s_60), .O(gate428inter3));
  inv1  gate971(.a(s_61), .O(gate428inter4));
  nand2 gate972(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate973(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate974(.a(G1048), .O(gate428inter7));
  inv1  gate975(.a(G1144), .O(gate428inter8));
  nand2 gate976(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate977(.a(s_61), .b(gate428inter3), .O(gate428inter10));
  nor2  gate978(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate979(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate980(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate883(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate884(.a(gate430inter0), .b(s_48), .O(gate430inter1));
  and2  gate885(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate886(.a(s_48), .O(gate430inter3));
  inv1  gate887(.a(s_49), .O(gate430inter4));
  nand2 gate888(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate889(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate890(.a(G1051), .O(gate430inter7));
  inv1  gate891(.a(G1147), .O(gate430inter8));
  nand2 gate892(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate893(.a(s_49), .b(gate430inter3), .O(gate430inter10));
  nor2  gate894(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate895(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate896(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate715(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate716(.a(gate433inter0), .b(s_24), .O(gate433inter1));
  and2  gate717(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate718(.a(s_24), .O(gate433inter3));
  inv1  gate719(.a(s_25), .O(gate433inter4));
  nand2 gate720(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate721(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate722(.a(G8), .O(gate433inter7));
  inv1  gate723(.a(G1153), .O(gate433inter8));
  nand2 gate724(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate725(.a(s_25), .b(gate433inter3), .O(gate433inter10));
  nor2  gate726(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate727(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate728(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1275(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1276(.a(gate438inter0), .b(s_104), .O(gate438inter1));
  and2  gate1277(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1278(.a(s_104), .O(gate438inter3));
  inv1  gate1279(.a(s_105), .O(gate438inter4));
  nand2 gate1280(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1281(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1282(.a(G1063), .O(gate438inter7));
  inv1  gate1283(.a(G1159), .O(gate438inter8));
  nand2 gate1284(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1285(.a(s_105), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1286(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1287(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1288(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate743(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate744(.a(gate441inter0), .b(s_28), .O(gate441inter1));
  and2  gate745(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate746(.a(s_28), .O(gate441inter3));
  inv1  gate747(.a(s_29), .O(gate441inter4));
  nand2 gate748(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate749(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate750(.a(G12), .O(gate441inter7));
  inv1  gate751(.a(G1165), .O(gate441inter8));
  nand2 gate752(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate753(.a(s_29), .b(gate441inter3), .O(gate441inter10));
  nor2  gate754(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate755(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate756(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate827(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate828(.a(gate449inter0), .b(s_40), .O(gate449inter1));
  and2  gate829(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate830(.a(s_40), .O(gate449inter3));
  inv1  gate831(.a(s_41), .O(gate449inter4));
  nand2 gate832(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate833(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate834(.a(G16), .O(gate449inter7));
  inv1  gate835(.a(G1177), .O(gate449inter8));
  nand2 gate836(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate837(.a(s_41), .b(gate449inter3), .O(gate449inter10));
  nor2  gate838(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate839(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate840(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate771(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate772(.a(gate450inter0), .b(s_32), .O(gate450inter1));
  and2  gate773(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate774(.a(s_32), .O(gate450inter3));
  inv1  gate775(.a(s_33), .O(gate450inter4));
  nand2 gate776(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate777(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate778(.a(G1081), .O(gate450inter7));
  inv1  gate779(.a(G1177), .O(gate450inter8));
  nand2 gate780(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate781(.a(s_33), .b(gate450inter3), .O(gate450inter10));
  nor2  gate782(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate783(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate784(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate603(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate604(.a(gate452inter0), .b(s_8), .O(gate452inter1));
  and2  gate605(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate606(.a(s_8), .O(gate452inter3));
  inv1  gate607(.a(s_9), .O(gate452inter4));
  nand2 gate608(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate609(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate610(.a(G1084), .O(gate452inter7));
  inv1  gate611(.a(G1180), .O(gate452inter8));
  nand2 gate612(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate613(.a(s_9), .b(gate452inter3), .O(gate452inter10));
  nor2  gate614(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate615(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate616(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1177(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1178(.a(gate455inter0), .b(s_90), .O(gate455inter1));
  and2  gate1179(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1180(.a(s_90), .O(gate455inter3));
  inv1  gate1181(.a(s_91), .O(gate455inter4));
  nand2 gate1182(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1183(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1184(.a(G19), .O(gate455inter7));
  inv1  gate1185(.a(G1186), .O(gate455inter8));
  nand2 gate1186(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1187(.a(s_91), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1188(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1189(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1190(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1975(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1976(.a(gate456inter0), .b(s_204), .O(gate456inter1));
  and2  gate1977(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1978(.a(s_204), .O(gate456inter3));
  inv1  gate1979(.a(s_205), .O(gate456inter4));
  nand2 gate1980(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1981(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1982(.a(G1090), .O(gate456inter7));
  inv1  gate1983(.a(G1186), .O(gate456inter8));
  nand2 gate1984(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1985(.a(s_205), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1986(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1987(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1988(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2031(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2032(.a(gate458inter0), .b(s_212), .O(gate458inter1));
  and2  gate2033(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2034(.a(s_212), .O(gate458inter3));
  inv1  gate2035(.a(s_213), .O(gate458inter4));
  nand2 gate2036(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2037(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2038(.a(G1093), .O(gate458inter7));
  inv1  gate2039(.a(G1189), .O(gate458inter8));
  nand2 gate2040(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2041(.a(s_213), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2042(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2043(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2044(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate855(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate856(.a(gate462inter0), .b(s_44), .O(gate462inter1));
  and2  gate857(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate858(.a(s_44), .O(gate462inter3));
  inv1  gate859(.a(s_45), .O(gate462inter4));
  nand2 gate860(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate861(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate862(.a(G1099), .O(gate462inter7));
  inv1  gate863(.a(G1195), .O(gate462inter8));
  nand2 gate864(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate865(.a(s_45), .b(gate462inter3), .O(gate462inter10));
  nor2  gate866(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate867(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate868(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2143(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2144(.a(gate463inter0), .b(s_228), .O(gate463inter1));
  and2  gate2145(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2146(.a(s_228), .O(gate463inter3));
  inv1  gate2147(.a(s_229), .O(gate463inter4));
  nand2 gate2148(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2149(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2150(.a(G23), .O(gate463inter7));
  inv1  gate2151(.a(G1198), .O(gate463inter8));
  nand2 gate2152(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2153(.a(s_229), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2154(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2155(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2156(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate757(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate758(.a(gate467inter0), .b(s_30), .O(gate467inter1));
  and2  gate759(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate760(.a(s_30), .O(gate467inter3));
  inv1  gate761(.a(s_31), .O(gate467inter4));
  nand2 gate762(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate763(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate764(.a(G25), .O(gate467inter7));
  inv1  gate765(.a(G1204), .O(gate467inter8));
  nand2 gate766(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate767(.a(s_31), .b(gate467inter3), .O(gate467inter10));
  nor2  gate768(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate769(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate770(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1331(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1332(.a(gate469inter0), .b(s_112), .O(gate469inter1));
  and2  gate1333(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1334(.a(s_112), .O(gate469inter3));
  inv1  gate1335(.a(s_113), .O(gate469inter4));
  nand2 gate1336(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1337(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1338(.a(G26), .O(gate469inter7));
  inv1  gate1339(.a(G1207), .O(gate469inter8));
  nand2 gate1340(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1341(.a(s_113), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1342(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1343(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1344(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate813(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate814(.a(gate470inter0), .b(s_38), .O(gate470inter1));
  and2  gate815(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate816(.a(s_38), .O(gate470inter3));
  inv1  gate817(.a(s_39), .O(gate470inter4));
  nand2 gate818(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate819(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate820(.a(G1111), .O(gate470inter7));
  inv1  gate821(.a(G1207), .O(gate470inter8));
  nand2 gate822(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate823(.a(s_39), .b(gate470inter3), .O(gate470inter10));
  nor2  gate824(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate825(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate826(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1345(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1346(.a(gate471inter0), .b(s_114), .O(gate471inter1));
  and2  gate1347(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1348(.a(s_114), .O(gate471inter3));
  inv1  gate1349(.a(s_115), .O(gate471inter4));
  nand2 gate1350(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1351(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1352(.a(G27), .O(gate471inter7));
  inv1  gate1353(.a(G1210), .O(gate471inter8));
  nand2 gate1354(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1355(.a(s_115), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1356(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1357(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1358(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate617(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate618(.a(gate477inter0), .b(s_10), .O(gate477inter1));
  and2  gate619(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate620(.a(s_10), .O(gate477inter3));
  inv1  gate621(.a(s_11), .O(gate477inter4));
  nand2 gate622(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate623(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate624(.a(G30), .O(gate477inter7));
  inv1  gate625(.a(G1219), .O(gate477inter8));
  nand2 gate626(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate627(.a(s_11), .b(gate477inter3), .O(gate477inter10));
  nor2  gate628(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate629(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate630(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate785(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate786(.a(gate479inter0), .b(s_34), .O(gate479inter1));
  and2  gate787(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate788(.a(s_34), .O(gate479inter3));
  inv1  gate789(.a(s_35), .O(gate479inter4));
  nand2 gate790(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate791(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate792(.a(G31), .O(gate479inter7));
  inv1  gate793(.a(G1222), .O(gate479inter8));
  nand2 gate794(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate795(.a(s_35), .b(gate479inter3), .O(gate479inter10));
  nor2  gate796(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate797(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate798(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1681(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1682(.a(gate481inter0), .b(s_162), .O(gate481inter1));
  and2  gate1683(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1684(.a(s_162), .O(gate481inter3));
  inv1  gate1685(.a(s_163), .O(gate481inter4));
  nand2 gate1686(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1687(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1688(.a(G32), .O(gate481inter7));
  inv1  gate1689(.a(G1225), .O(gate481inter8));
  nand2 gate1690(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1691(.a(s_163), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1692(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1693(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1694(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1121(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1122(.a(gate491inter0), .b(s_82), .O(gate491inter1));
  and2  gate1123(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1124(.a(s_82), .O(gate491inter3));
  inv1  gate1125(.a(s_83), .O(gate491inter4));
  nand2 gate1126(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1127(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1128(.a(G1244), .O(gate491inter7));
  inv1  gate1129(.a(G1245), .O(gate491inter8));
  nand2 gate1130(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1131(.a(s_83), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1132(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1133(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1134(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1583(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1584(.a(gate493inter0), .b(s_148), .O(gate493inter1));
  and2  gate1585(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1586(.a(s_148), .O(gate493inter3));
  inv1  gate1587(.a(s_149), .O(gate493inter4));
  nand2 gate1588(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1589(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1590(.a(G1248), .O(gate493inter7));
  inv1  gate1591(.a(G1249), .O(gate493inter8));
  nand2 gate1592(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1593(.a(s_149), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1594(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1595(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1596(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate645(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate646(.a(gate501inter0), .b(s_14), .O(gate501inter1));
  and2  gate647(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate648(.a(s_14), .O(gate501inter3));
  inv1  gate649(.a(s_15), .O(gate501inter4));
  nand2 gate650(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate651(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate652(.a(G1264), .O(gate501inter7));
  inv1  gate653(.a(G1265), .O(gate501inter8));
  nand2 gate654(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate655(.a(s_15), .b(gate501inter3), .O(gate501inter10));
  nor2  gate656(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate657(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate658(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1667(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1668(.a(gate502inter0), .b(s_160), .O(gate502inter1));
  and2  gate1669(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1670(.a(s_160), .O(gate502inter3));
  inv1  gate1671(.a(s_161), .O(gate502inter4));
  nand2 gate1672(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1673(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1674(.a(G1266), .O(gate502inter7));
  inv1  gate1675(.a(G1267), .O(gate502inter8));
  nand2 gate1676(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1677(.a(s_161), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1678(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1679(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1680(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate1863(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1864(.a(gate503inter0), .b(s_188), .O(gate503inter1));
  and2  gate1865(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1866(.a(s_188), .O(gate503inter3));
  inv1  gate1867(.a(s_189), .O(gate503inter4));
  nand2 gate1868(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1869(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1870(.a(G1268), .O(gate503inter7));
  inv1  gate1871(.a(G1269), .O(gate503inter8));
  nand2 gate1872(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1873(.a(s_189), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1874(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1875(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1876(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1597(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1598(.a(gate512inter0), .b(s_150), .O(gate512inter1));
  and2  gate1599(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1600(.a(s_150), .O(gate512inter3));
  inv1  gate1601(.a(s_151), .O(gate512inter4));
  nand2 gate1602(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1603(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1604(.a(G1286), .O(gate512inter7));
  inv1  gate1605(.a(G1287), .O(gate512inter8));
  nand2 gate1606(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1607(.a(s_151), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1608(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1609(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1610(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate673(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate674(.a(gate514inter0), .b(s_18), .O(gate514inter1));
  and2  gate675(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate676(.a(s_18), .O(gate514inter3));
  inv1  gate677(.a(s_19), .O(gate514inter4));
  nand2 gate678(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate679(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate680(.a(G1290), .O(gate514inter7));
  inv1  gate681(.a(G1291), .O(gate514inter8));
  nand2 gate682(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate683(.a(s_19), .b(gate514inter3), .O(gate514inter10));
  nor2  gate684(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate685(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate686(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule