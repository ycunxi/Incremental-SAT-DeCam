module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);

input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
input s_112,s_113;//RE__ALLOW(00,01,10,11);
input s_114,s_115;//RE__ALLOW(00,01,10,11);
input s_116,s_117;//RE__ALLOW(00,01,10,11);
input s_118,s_119;//RE__ALLOW(00,01,10,11);
input s_120,s_121;//RE__ALLOW(00,01,10,11);
input s_122,s_123;//RE__ALLOW(00,01,10,11);
input s_124,s_125;//RE__ALLOW(00,01,10,11);
input s_126,s_127;//RE__ALLOW(00,01,10,11);
input s_128,s_129;//RE__ALLOW(00,01,10,11);
input s_130,s_131;//RE__ALLOW(00,01,10,11);
input s_132,s_133;//RE__ALLOW(00,01,10,11);
input s_134,s_135;//RE__ALLOW(00,01,10,11);
input s_136,s_137;//RE__ALLOW(00,01,10,11);
input s_138,s_139;//RE__ALLOW(00,01,10,11);
input s_140,s_141;//RE__ALLOW(00,01,10,11);
input s_142,s_143;//RE__ALLOW(00,01,10,11);
input s_144,s_145;//RE__ALLOW(00,01,10,11);
input s_146,s_147;//RE__ALLOW(00,01,10,11);
input s_148,s_149;//RE__ALLOW(00,01,10,11);
input s_150,s_151;//RE__ALLOW(00,01,10,11);
input s_152,s_153;//RE__ALLOW(00,01,10,11);
input s_154,s_155;//RE__ALLOW(00,01,10,11);
input s_156,s_157;//RE__ALLOW(00,01,10,11);
input s_158,s_159;//RE__ALLOW(00,01,10,11);
input s_160,s_161;//RE__ALLOW(00,01,10,11);
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;

  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12;



and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1625(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1626(.a(gate9inter0), .b(s_154), .O(gate9inter1));
  and2  gate1627(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1628(.a(s_154), .O(gate9inter3));
  inv1  gate1629(.a(s_155), .O(gate9inter4));
  nand2 gate1630(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1631(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1632(.a(G1), .O(gate9inter7));
  inv1  gate1633(.a(G2), .O(gate9inter8));
  nand2 gate1634(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1635(.a(s_155), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1636(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1637(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1638(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1121(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1122(.a(gate17inter0), .b(s_82), .O(gate17inter1));
  and2  gate1123(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1124(.a(s_82), .O(gate17inter3));
  inv1  gate1125(.a(s_83), .O(gate17inter4));
  nand2 gate1126(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1127(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1128(.a(G17), .O(gate17inter7));
  inv1  gate1129(.a(G18), .O(gate17inter8));
  nand2 gate1130(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1131(.a(s_83), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1132(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1133(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1134(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate743(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate744(.a(gate26inter0), .b(s_28), .O(gate26inter1));
  and2  gate745(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate746(.a(s_28), .O(gate26inter3));
  inv1  gate747(.a(s_29), .O(gate26inter4));
  nand2 gate748(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate749(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate750(.a(G9), .O(gate26inter7));
  inv1  gate751(.a(G13), .O(gate26inter8));
  nand2 gate752(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate753(.a(s_29), .b(gate26inter3), .O(gate26inter10));
  nor2  gate754(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate755(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate756(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1359(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1360(.a(gate39inter0), .b(s_116), .O(gate39inter1));
  and2  gate1361(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1362(.a(s_116), .O(gate39inter3));
  inv1  gate1363(.a(s_117), .O(gate39inter4));
  nand2 gate1364(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1365(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1366(.a(G20), .O(gate39inter7));
  inv1  gate1367(.a(G24), .O(gate39inter8));
  nand2 gate1368(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1369(.a(s_117), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1370(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1371(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1372(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1429(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1430(.a(gate40inter0), .b(s_126), .O(gate40inter1));
  and2  gate1431(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1432(.a(s_126), .O(gate40inter3));
  inv1  gate1433(.a(s_127), .O(gate40inter4));
  nand2 gate1434(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1435(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1436(.a(G28), .O(gate40inter7));
  inv1  gate1437(.a(G32), .O(gate40inter8));
  nand2 gate1438(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1439(.a(s_127), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1440(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1441(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1442(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1289(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1290(.a(gate49inter0), .b(s_106), .O(gate49inter1));
  and2  gate1291(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1292(.a(s_106), .O(gate49inter3));
  inv1  gate1293(.a(s_107), .O(gate49inter4));
  nand2 gate1294(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1295(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1296(.a(G9), .O(gate49inter7));
  inv1  gate1297(.a(G278), .O(gate49inter8));
  nand2 gate1298(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1299(.a(s_107), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1300(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1301(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1302(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate925(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate926(.a(gate58inter0), .b(s_54), .O(gate58inter1));
  and2  gate927(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate928(.a(s_54), .O(gate58inter3));
  inv1  gate929(.a(s_55), .O(gate58inter4));
  nand2 gate930(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate931(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate932(.a(G18), .O(gate58inter7));
  inv1  gate933(.a(G290), .O(gate58inter8));
  nand2 gate934(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate935(.a(s_55), .b(gate58inter3), .O(gate58inter10));
  nor2  gate936(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate937(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate938(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1037(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1038(.a(gate66inter0), .b(s_70), .O(gate66inter1));
  and2  gate1039(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1040(.a(s_70), .O(gate66inter3));
  inv1  gate1041(.a(s_71), .O(gate66inter4));
  nand2 gate1042(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1043(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1044(.a(G26), .O(gate66inter7));
  inv1  gate1045(.a(G302), .O(gate66inter8));
  nand2 gate1046(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1047(.a(s_71), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1048(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1049(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1050(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1611(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1612(.a(gate70inter0), .b(s_152), .O(gate70inter1));
  and2  gate1613(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1614(.a(s_152), .O(gate70inter3));
  inv1  gate1615(.a(s_153), .O(gate70inter4));
  nand2 gate1616(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1617(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1618(.a(G30), .O(gate70inter7));
  inv1  gate1619(.a(G308), .O(gate70inter8));
  nand2 gate1620(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1621(.a(s_153), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1622(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1623(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1624(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate575(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate576(.a(gate74inter0), .b(s_4), .O(gate74inter1));
  and2  gate577(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate578(.a(s_4), .O(gate74inter3));
  inv1  gate579(.a(s_5), .O(gate74inter4));
  nand2 gate580(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate581(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate582(.a(G5), .O(gate74inter7));
  inv1  gate583(.a(G314), .O(gate74inter8));
  nand2 gate584(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate585(.a(s_5), .b(gate74inter3), .O(gate74inter10));
  nor2  gate586(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate587(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate588(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1555(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1556(.a(gate76inter0), .b(s_144), .O(gate76inter1));
  and2  gate1557(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1558(.a(s_144), .O(gate76inter3));
  inv1  gate1559(.a(s_145), .O(gate76inter4));
  nand2 gate1560(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1561(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1562(.a(G13), .O(gate76inter7));
  inv1  gate1563(.a(G317), .O(gate76inter8));
  nand2 gate1564(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1565(.a(s_145), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1566(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1567(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1568(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1639(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1640(.a(gate92inter0), .b(s_156), .O(gate92inter1));
  and2  gate1641(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1642(.a(s_156), .O(gate92inter3));
  inv1  gate1643(.a(s_157), .O(gate92inter4));
  nand2 gate1644(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1645(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1646(.a(G29), .O(gate92inter7));
  inv1  gate1647(.a(G341), .O(gate92inter8));
  nand2 gate1648(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1649(.a(s_157), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1650(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1651(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1652(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1107(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1108(.a(gate93inter0), .b(s_80), .O(gate93inter1));
  and2  gate1109(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1110(.a(s_80), .O(gate93inter3));
  inv1  gate1111(.a(s_81), .O(gate93inter4));
  nand2 gate1112(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1113(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1114(.a(G18), .O(gate93inter7));
  inv1  gate1115(.a(G344), .O(gate93inter8));
  nand2 gate1116(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1117(.a(s_81), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1118(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1119(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1120(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate673(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate674(.a(gate99inter0), .b(s_18), .O(gate99inter1));
  and2  gate675(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate676(.a(s_18), .O(gate99inter3));
  inv1  gate677(.a(s_19), .O(gate99inter4));
  nand2 gate678(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate679(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate680(.a(G27), .O(gate99inter7));
  inv1  gate681(.a(G353), .O(gate99inter8));
  nand2 gate682(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate683(.a(s_19), .b(gate99inter3), .O(gate99inter10));
  nor2  gate684(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate685(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate686(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1135(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1136(.a(gate106inter0), .b(s_84), .O(gate106inter1));
  and2  gate1137(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1138(.a(s_84), .O(gate106inter3));
  inv1  gate1139(.a(s_85), .O(gate106inter4));
  nand2 gate1140(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1141(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1142(.a(G364), .O(gate106inter7));
  inv1  gate1143(.a(G365), .O(gate106inter8));
  nand2 gate1144(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1145(.a(s_85), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1146(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1147(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1148(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate799(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate800(.a(gate108inter0), .b(s_36), .O(gate108inter1));
  and2  gate801(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate802(.a(s_36), .O(gate108inter3));
  inv1  gate803(.a(s_37), .O(gate108inter4));
  nand2 gate804(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate805(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate806(.a(G368), .O(gate108inter7));
  inv1  gate807(.a(G369), .O(gate108inter8));
  nand2 gate808(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate809(.a(s_37), .b(gate108inter3), .O(gate108inter10));
  nor2  gate810(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate811(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate812(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1317(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1318(.a(gate115inter0), .b(s_110), .O(gate115inter1));
  and2  gate1319(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1320(.a(s_110), .O(gate115inter3));
  inv1  gate1321(.a(s_111), .O(gate115inter4));
  nand2 gate1322(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1323(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1324(.a(G382), .O(gate115inter7));
  inv1  gate1325(.a(G383), .O(gate115inter8));
  nand2 gate1326(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1327(.a(s_111), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1328(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1329(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1330(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate981(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate982(.a(gate117inter0), .b(s_62), .O(gate117inter1));
  and2  gate983(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate984(.a(s_62), .O(gate117inter3));
  inv1  gate985(.a(s_63), .O(gate117inter4));
  nand2 gate986(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate987(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate988(.a(G386), .O(gate117inter7));
  inv1  gate989(.a(G387), .O(gate117inter8));
  nand2 gate990(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate991(.a(s_63), .b(gate117inter3), .O(gate117inter10));
  nor2  gate992(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate993(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate994(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1485(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1486(.a(gate120inter0), .b(s_134), .O(gate120inter1));
  and2  gate1487(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1488(.a(s_134), .O(gate120inter3));
  inv1  gate1489(.a(s_135), .O(gate120inter4));
  nand2 gate1490(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1491(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1492(.a(G392), .O(gate120inter7));
  inv1  gate1493(.a(G393), .O(gate120inter8));
  nand2 gate1494(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1495(.a(s_135), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1496(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1497(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1498(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate631(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate632(.a(gate123inter0), .b(s_12), .O(gate123inter1));
  and2  gate633(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate634(.a(s_12), .O(gate123inter3));
  inv1  gate635(.a(s_13), .O(gate123inter4));
  nand2 gate636(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate637(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate638(.a(G398), .O(gate123inter7));
  inv1  gate639(.a(G399), .O(gate123inter8));
  nand2 gate640(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate641(.a(s_13), .b(gate123inter3), .O(gate123inter10));
  nor2  gate642(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate643(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate644(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1233(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1234(.a(gate130inter0), .b(s_98), .O(gate130inter1));
  and2  gate1235(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1236(.a(s_98), .O(gate130inter3));
  inv1  gate1237(.a(s_99), .O(gate130inter4));
  nand2 gate1238(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1239(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1240(.a(G412), .O(gate130inter7));
  inv1  gate1241(.a(G413), .O(gate130inter8));
  nand2 gate1242(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1243(.a(s_99), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1244(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1245(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1246(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate715(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate716(.a(gate138inter0), .b(s_24), .O(gate138inter1));
  and2  gate717(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate718(.a(s_24), .O(gate138inter3));
  inv1  gate719(.a(s_25), .O(gate138inter4));
  nand2 gate720(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate721(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate722(.a(G432), .O(gate138inter7));
  inv1  gate723(.a(G435), .O(gate138inter8));
  nand2 gate724(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate725(.a(s_25), .b(gate138inter3), .O(gate138inter10));
  nor2  gate726(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate727(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate728(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate757(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate758(.a(gate157inter0), .b(s_30), .O(gate157inter1));
  and2  gate759(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate760(.a(s_30), .O(gate157inter3));
  inv1  gate761(.a(s_31), .O(gate157inter4));
  nand2 gate762(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate763(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate764(.a(G438), .O(gate157inter7));
  inv1  gate765(.a(G528), .O(gate157inter8));
  nand2 gate766(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate767(.a(s_31), .b(gate157inter3), .O(gate157inter10));
  nor2  gate768(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate769(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate770(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1303(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1304(.a(gate160inter0), .b(s_108), .O(gate160inter1));
  and2  gate1305(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1306(.a(s_108), .O(gate160inter3));
  inv1  gate1307(.a(s_109), .O(gate160inter4));
  nand2 gate1308(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1309(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1310(.a(G447), .O(gate160inter7));
  inv1  gate1311(.a(G531), .O(gate160inter8));
  nand2 gate1312(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1313(.a(s_109), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1314(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1315(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1316(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1261(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1262(.a(gate163inter0), .b(s_102), .O(gate163inter1));
  and2  gate1263(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1264(.a(s_102), .O(gate163inter3));
  inv1  gate1265(.a(s_103), .O(gate163inter4));
  nand2 gate1266(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1267(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1268(.a(G456), .O(gate163inter7));
  inv1  gate1269(.a(G537), .O(gate163inter8));
  nand2 gate1270(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1271(.a(s_103), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1272(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1273(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1274(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1093(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1094(.a(gate171inter0), .b(s_78), .O(gate171inter1));
  and2  gate1095(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1096(.a(s_78), .O(gate171inter3));
  inv1  gate1097(.a(s_79), .O(gate171inter4));
  nand2 gate1098(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1099(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1100(.a(G480), .O(gate171inter7));
  inv1  gate1101(.a(G549), .O(gate171inter8));
  nand2 gate1102(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1103(.a(s_79), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1104(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1105(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1106(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate701(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate702(.a(gate173inter0), .b(s_22), .O(gate173inter1));
  and2  gate703(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate704(.a(s_22), .O(gate173inter3));
  inv1  gate705(.a(s_23), .O(gate173inter4));
  nand2 gate706(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate707(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate708(.a(G486), .O(gate173inter7));
  inv1  gate709(.a(G552), .O(gate173inter8));
  nand2 gate710(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate711(.a(s_23), .b(gate173inter3), .O(gate173inter10));
  nor2  gate712(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate713(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate714(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1569(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1570(.a(gate178inter0), .b(s_146), .O(gate178inter1));
  and2  gate1571(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1572(.a(s_146), .O(gate178inter3));
  inv1  gate1573(.a(s_147), .O(gate178inter4));
  nand2 gate1574(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1575(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1576(.a(G501), .O(gate178inter7));
  inv1  gate1577(.a(G558), .O(gate178inter8));
  nand2 gate1578(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1579(.a(s_147), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1580(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1581(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1582(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate729(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate730(.a(gate180inter0), .b(s_26), .O(gate180inter1));
  and2  gate731(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate732(.a(s_26), .O(gate180inter3));
  inv1  gate733(.a(s_27), .O(gate180inter4));
  nand2 gate734(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate735(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate736(.a(G507), .O(gate180inter7));
  inv1  gate737(.a(G561), .O(gate180inter8));
  nand2 gate738(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate739(.a(s_27), .b(gate180inter3), .O(gate180inter10));
  nor2  gate740(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate741(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate742(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate771(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate772(.a(gate183inter0), .b(s_32), .O(gate183inter1));
  and2  gate773(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate774(.a(s_32), .O(gate183inter3));
  inv1  gate775(.a(s_33), .O(gate183inter4));
  nand2 gate776(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate777(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate778(.a(G516), .O(gate183inter7));
  inv1  gate779(.a(G567), .O(gate183inter8));
  nand2 gate780(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate781(.a(s_33), .b(gate183inter3), .O(gate183inter10));
  nor2  gate782(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate783(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate784(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate869(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate870(.a(gate186inter0), .b(s_46), .O(gate186inter1));
  and2  gate871(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate872(.a(s_46), .O(gate186inter3));
  inv1  gate873(.a(s_47), .O(gate186inter4));
  nand2 gate874(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate875(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate876(.a(G572), .O(gate186inter7));
  inv1  gate877(.a(G573), .O(gate186inter8));
  nand2 gate878(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate879(.a(s_47), .b(gate186inter3), .O(gate186inter10));
  nor2  gate880(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate881(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate882(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate1219(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1220(.a(gate194inter0), .b(s_96), .O(gate194inter1));
  and2  gate1221(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1222(.a(s_96), .O(gate194inter3));
  inv1  gate1223(.a(s_97), .O(gate194inter4));
  nand2 gate1224(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1225(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1226(.a(G588), .O(gate194inter7));
  inv1  gate1227(.a(G589), .O(gate194inter8));
  nand2 gate1228(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1229(.a(s_97), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1230(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1231(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1232(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1457(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1458(.a(gate195inter0), .b(s_130), .O(gate195inter1));
  and2  gate1459(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1460(.a(s_130), .O(gate195inter3));
  inv1  gate1461(.a(s_131), .O(gate195inter4));
  nand2 gate1462(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1463(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1464(.a(G590), .O(gate195inter7));
  inv1  gate1465(.a(G591), .O(gate195inter8));
  nand2 gate1466(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1467(.a(s_131), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1468(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1469(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1470(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1499(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1500(.a(gate203inter0), .b(s_136), .O(gate203inter1));
  and2  gate1501(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1502(.a(s_136), .O(gate203inter3));
  inv1  gate1503(.a(s_137), .O(gate203inter4));
  nand2 gate1504(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1505(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1506(.a(G602), .O(gate203inter7));
  inv1  gate1507(.a(G612), .O(gate203inter8));
  nand2 gate1508(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1509(.a(s_137), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1510(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1511(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1512(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1079(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1080(.a(gate205inter0), .b(s_76), .O(gate205inter1));
  and2  gate1081(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1082(.a(s_76), .O(gate205inter3));
  inv1  gate1083(.a(s_77), .O(gate205inter4));
  nand2 gate1084(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1085(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1086(.a(G622), .O(gate205inter7));
  inv1  gate1087(.a(G627), .O(gate205inter8));
  nand2 gate1088(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1089(.a(s_77), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1090(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1091(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1092(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1065(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1066(.a(gate212inter0), .b(s_74), .O(gate212inter1));
  and2  gate1067(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1068(.a(s_74), .O(gate212inter3));
  inv1  gate1069(.a(s_75), .O(gate212inter4));
  nand2 gate1070(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1071(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1072(.a(G617), .O(gate212inter7));
  inv1  gate1073(.a(G669), .O(gate212inter8));
  nand2 gate1074(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1075(.a(s_75), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1076(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1077(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1078(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1191(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1192(.a(gate215inter0), .b(s_92), .O(gate215inter1));
  and2  gate1193(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1194(.a(s_92), .O(gate215inter3));
  inv1  gate1195(.a(s_93), .O(gate215inter4));
  nand2 gate1196(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1197(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1198(.a(G607), .O(gate215inter7));
  inv1  gate1199(.a(G675), .O(gate215inter8));
  nand2 gate1200(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1201(.a(s_93), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1202(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1203(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1204(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate617(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate618(.a(gate223inter0), .b(s_10), .O(gate223inter1));
  and2  gate619(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate620(.a(s_10), .O(gate223inter3));
  inv1  gate621(.a(s_11), .O(gate223inter4));
  nand2 gate622(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate623(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate624(.a(G627), .O(gate223inter7));
  inv1  gate625(.a(G687), .O(gate223inter8));
  nand2 gate626(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate627(.a(s_11), .b(gate223inter3), .O(gate223inter10));
  nor2  gate628(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate629(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate630(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1653(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1654(.a(gate224inter0), .b(s_158), .O(gate224inter1));
  and2  gate1655(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1656(.a(s_158), .O(gate224inter3));
  inv1  gate1657(.a(s_159), .O(gate224inter4));
  nand2 gate1658(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1659(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1660(.a(G637), .O(gate224inter7));
  inv1  gate1661(.a(G687), .O(gate224inter8));
  nand2 gate1662(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1663(.a(s_159), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1664(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1665(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1666(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1149(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1150(.a(gate227inter0), .b(s_86), .O(gate227inter1));
  and2  gate1151(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1152(.a(s_86), .O(gate227inter3));
  inv1  gate1153(.a(s_87), .O(gate227inter4));
  nand2 gate1154(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1155(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1156(.a(G694), .O(gate227inter7));
  inv1  gate1157(.a(G695), .O(gate227inter8));
  nand2 gate1158(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1159(.a(s_87), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1160(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1161(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1162(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate645(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate646(.a(gate243inter0), .b(s_14), .O(gate243inter1));
  and2  gate647(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate648(.a(s_14), .O(gate243inter3));
  inv1  gate649(.a(s_15), .O(gate243inter4));
  nand2 gate650(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate651(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate652(.a(G245), .O(gate243inter7));
  inv1  gate653(.a(G733), .O(gate243inter8));
  nand2 gate654(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate655(.a(s_15), .b(gate243inter3), .O(gate243inter10));
  nor2  gate656(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate657(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate658(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1667(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1668(.a(gate248inter0), .b(s_160), .O(gate248inter1));
  and2  gate1669(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1670(.a(s_160), .O(gate248inter3));
  inv1  gate1671(.a(s_161), .O(gate248inter4));
  nand2 gate1672(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1673(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1674(.a(G727), .O(gate248inter7));
  inv1  gate1675(.a(G739), .O(gate248inter8));
  nand2 gate1676(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1677(.a(s_161), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1678(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1679(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1680(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1541(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1542(.a(gate264inter0), .b(s_142), .O(gate264inter1));
  and2  gate1543(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1544(.a(s_142), .O(gate264inter3));
  inv1  gate1545(.a(s_143), .O(gate264inter4));
  nand2 gate1546(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1547(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1548(.a(G768), .O(gate264inter7));
  inv1  gate1549(.a(G769), .O(gate264inter8));
  nand2 gate1550(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1551(.a(s_143), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1552(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1553(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1554(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1163(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1164(.a(gate271inter0), .b(s_88), .O(gate271inter1));
  and2  gate1165(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1166(.a(s_88), .O(gate271inter3));
  inv1  gate1167(.a(s_89), .O(gate271inter4));
  nand2 gate1168(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1169(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1170(.a(G660), .O(gate271inter7));
  inv1  gate1171(.a(G788), .O(gate271inter8));
  nand2 gate1172(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1173(.a(s_89), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1174(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1175(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1176(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1331(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1332(.a(gate274inter0), .b(s_112), .O(gate274inter1));
  and2  gate1333(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1334(.a(s_112), .O(gate274inter3));
  inv1  gate1335(.a(s_113), .O(gate274inter4));
  nand2 gate1336(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1337(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1338(.a(G770), .O(gate274inter7));
  inv1  gate1339(.a(G794), .O(gate274inter8));
  nand2 gate1340(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1341(.a(s_113), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1342(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1343(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1344(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1275(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1276(.a(gate276inter0), .b(s_104), .O(gate276inter1));
  and2  gate1277(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1278(.a(s_104), .O(gate276inter3));
  inv1  gate1279(.a(s_105), .O(gate276inter4));
  nand2 gate1280(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1281(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1282(.a(G773), .O(gate276inter7));
  inv1  gate1283(.a(G797), .O(gate276inter8));
  nand2 gate1284(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1285(.a(s_105), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1286(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1287(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1288(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1597(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1598(.a(gate284inter0), .b(s_150), .O(gate284inter1));
  and2  gate1599(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1600(.a(s_150), .O(gate284inter3));
  inv1  gate1601(.a(s_151), .O(gate284inter4));
  nand2 gate1602(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1603(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1604(.a(G785), .O(gate284inter7));
  inv1  gate1605(.a(G809), .O(gate284inter8));
  nand2 gate1606(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1607(.a(s_151), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1608(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1609(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1610(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate813(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate814(.a(gate286inter0), .b(s_38), .O(gate286inter1));
  and2  gate815(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate816(.a(s_38), .O(gate286inter3));
  inv1  gate817(.a(s_39), .O(gate286inter4));
  nand2 gate818(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate819(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate820(.a(G788), .O(gate286inter7));
  inv1  gate821(.a(G812), .O(gate286inter8));
  nand2 gate822(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate823(.a(s_39), .b(gate286inter3), .O(gate286inter10));
  nor2  gate824(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate825(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate826(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1583(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1584(.a(gate287inter0), .b(s_148), .O(gate287inter1));
  and2  gate1585(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1586(.a(s_148), .O(gate287inter3));
  inv1  gate1587(.a(s_149), .O(gate287inter4));
  nand2 gate1588(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1589(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1590(.a(G663), .O(gate287inter7));
  inv1  gate1591(.a(G815), .O(gate287inter8));
  nand2 gate1592(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1593(.a(s_149), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1594(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1595(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1596(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate953(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate954(.a(gate289inter0), .b(s_58), .O(gate289inter1));
  and2  gate955(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate956(.a(s_58), .O(gate289inter3));
  inv1  gate957(.a(s_59), .O(gate289inter4));
  nand2 gate958(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate959(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate960(.a(G818), .O(gate289inter7));
  inv1  gate961(.a(G819), .O(gate289inter8));
  nand2 gate962(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate963(.a(s_59), .b(gate289inter3), .O(gate289inter10));
  nor2  gate964(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate965(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate966(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate939(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate940(.a(gate290inter0), .b(s_56), .O(gate290inter1));
  and2  gate941(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate942(.a(s_56), .O(gate290inter3));
  inv1  gate943(.a(s_57), .O(gate290inter4));
  nand2 gate944(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate945(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate946(.a(G820), .O(gate290inter7));
  inv1  gate947(.a(G821), .O(gate290inter8));
  nand2 gate948(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate949(.a(s_57), .b(gate290inter3), .O(gate290inter10));
  nor2  gate950(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate951(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate952(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1415(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1416(.a(gate295inter0), .b(s_124), .O(gate295inter1));
  and2  gate1417(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1418(.a(s_124), .O(gate295inter3));
  inv1  gate1419(.a(s_125), .O(gate295inter4));
  nand2 gate1420(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1421(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1422(.a(G830), .O(gate295inter7));
  inv1  gate1423(.a(G831), .O(gate295inter8));
  nand2 gate1424(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1425(.a(s_125), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1426(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1427(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1428(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate589(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate590(.a(gate390inter0), .b(s_6), .O(gate390inter1));
  and2  gate591(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate592(.a(s_6), .O(gate390inter3));
  inv1  gate593(.a(s_7), .O(gate390inter4));
  nand2 gate594(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate595(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate596(.a(G4), .O(gate390inter7));
  inv1  gate597(.a(G1045), .O(gate390inter8));
  nand2 gate598(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate599(.a(s_7), .b(gate390inter3), .O(gate390inter10));
  nor2  gate600(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate601(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate602(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate561(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate562(.a(gate391inter0), .b(s_2), .O(gate391inter1));
  and2  gate563(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate564(.a(s_2), .O(gate391inter3));
  inv1  gate565(.a(s_3), .O(gate391inter4));
  nand2 gate566(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate567(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate568(.a(G5), .O(gate391inter7));
  inv1  gate569(.a(G1048), .O(gate391inter8));
  nand2 gate570(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate571(.a(s_3), .b(gate391inter3), .O(gate391inter10));
  nor2  gate572(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate573(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate574(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate827(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate828(.a(gate404inter0), .b(s_40), .O(gate404inter1));
  and2  gate829(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate830(.a(s_40), .O(gate404inter3));
  inv1  gate831(.a(s_41), .O(gate404inter4));
  nand2 gate832(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate833(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate834(.a(G18), .O(gate404inter7));
  inv1  gate835(.a(G1087), .O(gate404inter8));
  nand2 gate836(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate837(.a(s_41), .b(gate404inter3), .O(gate404inter10));
  nor2  gate838(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate839(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate840(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate841(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate842(.a(gate410inter0), .b(s_42), .O(gate410inter1));
  and2  gate843(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate844(.a(s_42), .O(gate410inter3));
  inv1  gate845(.a(s_43), .O(gate410inter4));
  nand2 gate846(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate847(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate848(.a(G24), .O(gate410inter7));
  inv1  gate849(.a(G1105), .O(gate410inter8));
  nand2 gate850(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate851(.a(s_43), .b(gate410inter3), .O(gate410inter10));
  nor2  gate852(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate853(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate854(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate855(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate856(.a(gate412inter0), .b(s_44), .O(gate412inter1));
  and2  gate857(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate858(.a(s_44), .O(gate412inter3));
  inv1  gate859(.a(s_45), .O(gate412inter4));
  nand2 gate860(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate861(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate862(.a(G26), .O(gate412inter7));
  inv1  gate863(.a(G1111), .O(gate412inter8));
  nand2 gate864(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate865(.a(s_45), .b(gate412inter3), .O(gate412inter10));
  nor2  gate866(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate867(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate868(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1345(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1346(.a(gate415inter0), .b(s_114), .O(gate415inter1));
  and2  gate1347(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1348(.a(s_114), .O(gate415inter3));
  inv1  gate1349(.a(s_115), .O(gate415inter4));
  nand2 gate1350(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1351(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1352(.a(G29), .O(gate415inter7));
  inv1  gate1353(.a(G1120), .O(gate415inter8));
  nand2 gate1354(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1355(.a(s_115), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1356(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1357(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1358(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1373(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1374(.a(gate423inter0), .b(s_118), .O(gate423inter1));
  and2  gate1375(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1376(.a(s_118), .O(gate423inter3));
  inv1  gate1377(.a(s_119), .O(gate423inter4));
  nand2 gate1378(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1379(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1380(.a(G3), .O(gate423inter7));
  inv1  gate1381(.a(G1138), .O(gate423inter8));
  nand2 gate1382(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1383(.a(s_119), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1384(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1385(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1386(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1023(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1024(.a(gate427inter0), .b(s_68), .O(gate427inter1));
  and2  gate1025(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1026(.a(s_68), .O(gate427inter3));
  inv1  gate1027(.a(s_69), .O(gate427inter4));
  nand2 gate1028(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1029(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1030(.a(G5), .O(gate427inter7));
  inv1  gate1031(.a(G1144), .O(gate427inter8));
  nand2 gate1032(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1033(.a(s_69), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1034(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1035(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1036(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1471(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1472(.a(gate431inter0), .b(s_132), .O(gate431inter1));
  and2  gate1473(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1474(.a(s_132), .O(gate431inter3));
  inv1  gate1475(.a(s_133), .O(gate431inter4));
  nand2 gate1476(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1477(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1478(.a(G7), .O(gate431inter7));
  inv1  gate1479(.a(G1150), .O(gate431inter8));
  nand2 gate1480(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1481(.a(s_133), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1482(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1483(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1484(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1051(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1052(.a(gate433inter0), .b(s_72), .O(gate433inter1));
  and2  gate1053(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1054(.a(s_72), .O(gate433inter3));
  inv1  gate1055(.a(s_73), .O(gate433inter4));
  nand2 gate1056(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1057(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1058(.a(G8), .O(gate433inter7));
  inv1  gate1059(.a(G1153), .O(gate433inter8));
  nand2 gate1060(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1061(.a(s_73), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1062(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1063(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1064(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate603(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate604(.a(gate434inter0), .b(s_8), .O(gate434inter1));
  and2  gate605(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate606(.a(s_8), .O(gate434inter3));
  inv1  gate607(.a(s_9), .O(gate434inter4));
  nand2 gate608(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate609(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate610(.a(G1057), .O(gate434inter7));
  inv1  gate611(.a(G1153), .O(gate434inter8));
  nand2 gate612(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate613(.a(s_9), .b(gate434inter3), .O(gate434inter10));
  nor2  gate614(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate615(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate616(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate547(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate548(.a(gate437inter0), .b(s_0), .O(gate437inter1));
  and2  gate549(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate550(.a(s_0), .O(gate437inter3));
  inv1  gate551(.a(s_1), .O(gate437inter4));
  nand2 gate552(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate553(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate554(.a(G10), .O(gate437inter7));
  inv1  gate555(.a(G1159), .O(gate437inter8));
  nand2 gate556(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate557(.a(s_1), .b(gate437inter3), .O(gate437inter10));
  nor2  gate558(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate559(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate560(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1527(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1528(.a(gate442inter0), .b(s_140), .O(gate442inter1));
  and2  gate1529(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1530(.a(s_140), .O(gate442inter3));
  inv1  gate1531(.a(s_141), .O(gate442inter4));
  nand2 gate1532(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1533(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1534(.a(G1069), .O(gate442inter7));
  inv1  gate1535(.a(G1165), .O(gate442inter8));
  nand2 gate1536(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1537(.a(s_141), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1538(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1539(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1540(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1177(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1178(.a(gate445inter0), .b(s_90), .O(gate445inter1));
  and2  gate1179(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1180(.a(s_90), .O(gate445inter3));
  inv1  gate1181(.a(s_91), .O(gate445inter4));
  nand2 gate1182(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1183(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1184(.a(G14), .O(gate445inter7));
  inv1  gate1185(.a(G1171), .O(gate445inter8));
  nand2 gate1186(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1187(.a(s_91), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1188(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1189(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1190(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate883(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate884(.a(gate448inter0), .b(s_48), .O(gate448inter1));
  and2  gate885(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate886(.a(s_48), .O(gate448inter3));
  inv1  gate887(.a(s_49), .O(gate448inter4));
  nand2 gate888(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate889(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate890(.a(G1078), .O(gate448inter7));
  inv1  gate891(.a(G1174), .O(gate448inter8));
  nand2 gate892(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate893(.a(s_49), .b(gate448inter3), .O(gate448inter10));
  nor2  gate894(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate895(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate896(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate659(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate660(.a(gate449inter0), .b(s_16), .O(gate449inter1));
  and2  gate661(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate662(.a(s_16), .O(gate449inter3));
  inv1  gate663(.a(s_17), .O(gate449inter4));
  nand2 gate664(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate665(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate666(.a(G16), .O(gate449inter7));
  inv1  gate667(.a(G1177), .O(gate449inter8));
  nand2 gate668(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate669(.a(s_17), .b(gate449inter3), .O(gate449inter10));
  nor2  gate670(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate671(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate672(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1387(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1388(.a(gate464inter0), .b(s_120), .O(gate464inter1));
  and2  gate1389(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1390(.a(s_120), .O(gate464inter3));
  inv1  gate1391(.a(s_121), .O(gate464inter4));
  nand2 gate1392(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1393(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1394(.a(G1102), .O(gate464inter7));
  inv1  gate1395(.a(G1198), .O(gate464inter8));
  nand2 gate1396(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1397(.a(s_121), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1398(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1399(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1400(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate897(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate898(.a(gate465inter0), .b(s_50), .O(gate465inter1));
  and2  gate899(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate900(.a(s_50), .O(gate465inter3));
  inv1  gate901(.a(s_51), .O(gate465inter4));
  nand2 gate902(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate903(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate904(.a(G24), .O(gate465inter7));
  inv1  gate905(.a(G1201), .O(gate465inter8));
  nand2 gate906(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate907(.a(s_51), .b(gate465inter3), .O(gate465inter10));
  nor2  gate908(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate909(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate910(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate995(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate996(.a(gate470inter0), .b(s_64), .O(gate470inter1));
  and2  gate997(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate998(.a(s_64), .O(gate470inter3));
  inv1  gate999(.a(s_65), .O(gate470inter4));
  nand2 gate1000(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1001(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1002(.a(G1111), .O(gate470inter7));
  inv1  gate1003(.a(G1207), .O(gate470inter8));
  nand2 gate1004(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1005(.a(s_65), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1006(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1007(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1008(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1205(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1206(.a(gate471inter0), .b(s_94), .O(gate471inter1));
  and2  gate1207(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1208(.a(s_94), .O(gate471inter3));
  inv1  gate1209(.a(s_95), .O(gate471inter4));
  nand2 gate1210(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1211(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1212(.a(G27), .O(gate471inter7));
  inv1  gate1213(.a(G1210), .O(gate471inter8));
  nand2 gate1214(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1215(.a(s_95), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1216(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1217(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1218(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1247(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1248(.a(gate476inter0), .b(s_100), .O(gate476inter1));
  and2  gate1249(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1250(.a(s_100), .O(gate476inter3));
  inv1  gate1251(.a(s_101), .O(gate476inter4));
  nand2 gate1252(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1253(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1254(.a(G1120), .O(gate476inter7));
  inv1  gate1255(.a(G1216), .O(gate476inter8));
  nand2 gate1256(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1257(.a(s_101), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1258(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1259(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1260(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1513(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1514(.a(gate478inter0), .b(s_138), .O(gate478inter1));
  and2  gate1515(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1516(.a(s_138), .O(gate478inter3));
  inv1  gate1517(.a(s_139), .O(gate478inter4));
  nand2 gate1518(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1519(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1520(.a(G1123), .O(gate478inter7));
  inv1  gate1521(.a(G1219), .O(gate478inter8));
  nand2 gate1522(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1523(.a(s_139), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1524(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1525(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1526(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate967(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate968(.a(gate479inter0), .b(s_60), .O(gate479inter1));
  and2  gate969(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate970(.a(s_60), .O(gate479inter3));
  inv1  gate971(.a(s_61), .O(gate479inter4));
  nand2 gate972(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate973(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate974(.a(G31), .O(gate479inter7));
  inv1  gate975(.a(G1222), .O(gate479inter8));
  nand2 gate976(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate977(.a(s_61), .b(gate479inter3), .O(gate479inter10));
  nor2  gate978(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate979(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate980(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate911(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate912(.a(gate481inter0), .b(s_52), .O(gate481inter1));
  and2  gate913(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate914(.a(s_52), .O(gate481inter3));
  inv1  gate915(.a(s_53), .O(gate481inter4));
  nand2 gate916(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate917(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate918(.a(G32), .O(gate481inter7));
  inv1  gate919(.a(G1225), .O(gate481inter8));
  nand2 gate920(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate921(.a(s_53), .b(gate481inter3), .O(gate481inter10));
  nor2  gate922(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate923(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate924(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate687(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate688(.a(gate487inter0), .b(s_20), .O(gate487inter1));
  and2  gate689(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate690(.a(s_20), .O(gate487inter3));
  inv1  gate691(.a(s_21), .O(gate487inter4));
  nand2 gate692(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate693(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate694(.a(G1236), .O(gate487inter7));
  inv1  gate695(.a(G1237), .O(gate487inter8));
  nand2 gate696(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate697(.a(s_21), .b(gate487inter3), .O(gate487inter10));
  nor2  gate698(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate699(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate700(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1401(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1402(.a(gate495inter0), .b(s_122), .O(gate495inter1));
  and2  gate1403(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1404(.a(s_122), .O(gate495inter3));
  inv1  gate1405(.a(s_123), .O(gate495inter4));
  nand2 gate1406(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1407(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1408(.a(G1252), .O(gate495inter7));
  inv1  gate1409(.a(G1253), .O(gate495inter8));
  nand2 gate1410(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1411(.a(s_123), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1412(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1413(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1414(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1009(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1010(.a(gate506inter0), .b(s_66), .O(gate506inter1));
  and2  gate1011(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1012(.a(s_66), .O(gate506inter3));
  inv1  gate1013(.a(s_67), .O(gate506inter4));
  nand2 gate1014(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1015(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1016(.a(G1274), .O(gate506inter7));
  inv1  gate1017(.a(G1275), .O(gate506inter8));
  nand2 gate1018(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1019(.a(s_67), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1020(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1021(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1022(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate1443(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate1444(.a(gate513inter0), .b(s_128), .O(gate513inter1));
  and2  gate1445(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate1446(.a(s_128), .O(gate513inter3));
  inv1  gate1447(.a(s_129), .O(gate513inter4));
  nand2 gate1448(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate1449(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate1450(.a(G1288), .O(gate513inter7));
  inv1  gate1451(.a(G1289), .O(gate513inter8));
  nand2 gate1452(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate1453(.a(s_129), .b(gate513inter3), .O(gate513inter10));
  nor2  gate1454(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate1455(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate1456(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate785(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate786(.a(gate514inter0), .b(s_34), .O(gate514inter1));
  and2  gate787(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate788(.a(s_34), .O(gate514inter3));
  inv1  gate789(.a(s_35), .O(gate514inter4));
  nand2 gate790(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate791(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate792(.a(G1290), .O(gate514inter7));
  inv1  gate793(.a(G1291), .O(gate514inter8));
  nand2 gate794(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate795(.a(s_35), .b(gate514inter3), .O(gate514inter10));
  nor2  gate796(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate797(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate798(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule