module c2670 (N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
              N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
              N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
              N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
              N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
              N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
              N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
              N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
              N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
              N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
              N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
              N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
              N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
              N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
              N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
              N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
              N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
              N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
              N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
              N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
              N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
              N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
              N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
              N216_I,N217_I,N218_I,N398,N400,N401,N419,N420,N456,N457,
              N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,
              N799,N805,N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,
              N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,
              N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,
              N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,
              N3803,N3804,N3809,N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,
              N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,
              N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,
              N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,
              N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,
              N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,
              N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,
              N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,
              N216_O,N217_O,N218_O);

input N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
      N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
      N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
      N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
      N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
      N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
      N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
      N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
      N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
      N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
      N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
      N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
      N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
      N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
      N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
      N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
      N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
      N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
      N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
      N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
      N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
      N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
      N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
      N216_I,N217_I,N218_I;//RE__PI;

input s_0,s_1;//RE__ALLOW(00,01,10,11);
input s_2,s_3;//RE__ALLOW(00,01,10,11);
input s_4,s_5;//RE__ALLOW(00,01,10,11);
input s_6,s_7;//RE__ALLOW(00,01,10,11);
input s_8,s_9;//RE__ALLOW(00,01,10,11);
input s_10,s_11;//RE__ALLOW(00,01,10,11);
input s_12,s_13;//RE__ALLOW(00,01,10,11);
input s_14,s_15;//RE__ALLOW(00,01,10,11);
input s_16,s_17;//RE__ALLOW(00,01,10,11);
input s_18,s_19;//RE__ALLOW(00,01,10,11);
input s_20,s_21;//RE__ALLOW(00,01,10,11);
input s_22,s_23;//RE__ALLOW(00,01,10,11);
input s_24,s_25;//RE__ALLOW(00,01,10,11);
input s_26,s_27;//RE__ALLOW(00,01,10,11);
input s_28,s_29;//RE__ALLOW(00,01,10,11);
input s_30,s_31;//RE__ALLOW(00,01,10,11);
input s_32,s_33;//RE__ALLOW(00,01,10,11);
input s_34,s_35;//RE__ALLOW(00,01,10,11);
input s_36,s_37;//RE__ALLOW(00,01,10,11);
input s_38,s_39;//RE__ALLOW(00,01,10,11);
input s_40,s_41;//RE__ALLOW(00,01,10,11);
input s_42,s_43;//RE__ALLOW(00,01,10,11);
input s_44,s_45;//RE__ALLOW(00,01,10,11);
input s_46,s_47;//RE__ALLOW(00,01,10,11);
input s_48,s_49;//RE__ALLOW(00,01,10,11);
input s_50,s_51;//RE__ALLOW(00,01,10,11);
input s_52,s_53;//RE__ALLOW(00,01,10,11);
input s_54,s_55;//RE__ALLOW(00,01,10,11);
input s_56,s_57;//RE__ALLOW(00,01,10,11);
input s_58,s_59;//RE__ALLOW(00,01,10,11);
input s_60,s_61;//RE__ALLOW(00,01,10,11);
input s_62,s_63;//RE__ALLOW(00,01,10,11);
input s_64,s_65;//RE__ALLOW(00,01,10,11);
input s_66,s_67;//RE__ALLOW(00,01,10,11);
input s_68,s_69;//RE__ALLOW(00,01,10,11);
input s_70,s_71;//RE__ALLOW(00,01,10,11);
input s_72,s_73;//RE__ALLOW(00,01,10,11);
input s_74,s_75;//RE__ALLOW(00,01,10,11);
input s_76,s_77;//RE__ALLOW(00,01,10,11);
input s_78,s_79;//RE__ALLOW(00,01,10,11);
input s_80,s_81;//RE__ALLOW(00,01,10,11);
input s_82,s_83;//RE__ALLOW(00,01,10,11);
input s_84,s_85;//RE__ALLOW(00,01,10,11);
input s_86,s_87;//RE__ALLOW(00,01,10,11);
input s_88,s_89;//RE__ALLOW(00,01,10,11);
input s_90,s_91;//RE__ALLOW(00,01,10,11);
input s_92,s_93;//RE__ALLOW(00,01,10,11);
input s_94,s_95;//RE__ALLOW(00,01,10,11);
input s_96,s_97;//RE__ALLOW(00,01,10,11);
input s_98,s_99;//RE__ALLOW(00,01,10,11);
input s_100,s_101;//RE__ALLOW(00,01,10,11);
input s_102,s_103;//RE__ALLOW(00,01,10,11);
input s_104,s_105;//RE__ALLOW(00,01,10,11);
input s_106,s_107;//RE__ALLOW(00,01,10,11);
input s_108,s_109;//RE__ALLOW(00,01,10,11);
input s_110,s_111;//RE__ALLOW(00,01,10,11);
output N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,
       N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,
       N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,
       N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,
       N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,
       N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,
       N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,
       N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,
       N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,
       N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,
       N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,
       N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,
       N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,
       N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O;

wire N405,N408,N425,N485,N486,N495,N496,N499,N500,N503,
     N506,N509,N521,N533,N537,N543,N544,N547,N550,N562,
     N574,N578,N582,N594,N606,N607,N608,N609,N610,N611,
     N612,N613,N625,N637,N643,N650,N651,N655,N659,N663,
     N667,N671,N675,N679,N683,N687,N693,N699,N705,N711,
     N715,N719,N723,N727,N730,N733,N734,N735,N738,N741,
     N744,N747,N750,N753,N756,N759,N762,N765,N768,N771,
     N774,N777,N780,N783,N786,N800,N900,N901,N902,N903,
     N904,N905,N998,N999,N1027,N1032,N1033,N1034,N1037,N1042,
     N1053,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1075,N1086,
     N1097,N1098,N1099,N1100,N1101,N1102,N1113,N1124,N1125,N1126,
     N1127,N1128,N1129,N1133,N1137,N1140,N1141,N1142,N1143,N1144,
     N1145,N1146,N1157,N1168,N1169,N1170,N1171,N1172,N1173,N1178,
     N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1195,N1200,N1205,
     N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1219,N1222,N1225,
     N1228,N1231,N1234,N1237,N1240,N1243,N1246,N1249,N1250,N1251,
     N1254,N1257,N1260,N1263,N1266,N1275,N1276,N1302,N1351,N1352,
     N1353,N1354,N1355,N1395,N1396,N1397,N1398,N1399,N1422,N1423,
     N1424,N1425,N1426,N1427,N1440,N1441,N1449,N1450,N1451,N1452,
     N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,
     N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
     N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,
     N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,
     N1493,N1494,N1495,N1496,N1499,N1502,N1506,N1510,N1513,N1516,
     N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
     N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
     N1549,N1550,N1551,N1552,N1553,N1557,N1561,N1564,N1565,N1566,
     N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,
     N1577,N1578,N1581,N1582,N1585,N1588,N1591,N1596,N1600,N1606,
     N1612,N1615,N1619,N1624,N1628,N1631,N1634,N1637,N1642,N1647,
     N1651,N1656,N1676,N1681,N1686,N1690,N1708,N1770,N1773,N1776,
     N1777,N1778,N1781,N1784,N1785,N1795,N1798,N1801,N1804,N1807,
     N1808,N1809,N1810,N1811,N1813,N1814,N1815,N1822,N1823,N1824,
     N1827,N1830,N1831,N1832,N1833,N1836,N1841,N1848,N1852,N1856,
     N1863,N1870,N1875,N1880,N1885,N1888,N1891,N1894,N1897,N1908,
     N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,
     N1919,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,
     N1939,N1940,N1941,N1942,N1945,N1948,N1951,N1954,N1957,N1960,
     N1963,N1966,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2040,
     N2041,N2042,N2043,N2046,N2049,N2052,N2055,N2058,N2061,N2064,
     N2067,N2070,N2073,N2076,N2079,N2095,N2098,N2101,N2104,N2107,
     N2110,N2113,N2119,N2120,N2125,N2126,N2127,N2128,N2135,N2141,
     N2144,N2147,N2150,N2153,N2154,N2155,N2156,N2157,N2158,N2171,
     N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2185,N2188,N2191,
     N2194,N2197,N2200,N2201,N2204,N2207,N2210,N2213,N2216,N2219,
     N2234,N2235,N2236,N2237,N2250,N2266,N2269,N2291,N2294,N2297,
     N2298,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,
     N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,
     N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,
     N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
     N2339,N2340,N2354,N2355,N2356,N2357,N2358,N2359,N2364,N2365,
     N2366,N2367,N2368,N2372,N2373,N2374,N2375,N2376,N2377,N2382,
     N2386,N2391,N2395,N2400,N2403,N2406,N2407,N2408,N2409,N2410,
     N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2421,N2425,N2428,
     N2429,N2430,N2431,N2432,N2433,N2434,N2437,N2440,N2443,N2446,
     N2449,N2452,N2453,N2454,N2457,N2460,N2463,N2466,N2469,N2472,
     N2475,N2478,N2481,N2484,N2487,N2490,N2493,N2503,N2504,N2510,
     N2511,N2521,N2528,N2531,N2534,N2537,N2540,N2544,N2545,N2546,
     N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2563,N2564,N2565,
     N2566,N2567,N2568,N2579,N2603,N2607,N2608,N2609,N2610,N2611,
     N2612,N2613,N2617,N2618,N2619,N2620,N2621,N2624,N2628,N2629,
     N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2638,N2645,N2646,
     N2652,N2655,N2656,N2659,N2663,N2664,N2665,N2666,N2667,N2668,
     N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,
     N2679,N2680,N2681,N2684,N2687,N2690,N2693,N2694,N2695,N2696,
     N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2706,N2707,N2708,
     N2709,N2710,N2719,N2720,N2726,N2729,N2738,N2743,N2747,N2748,
     N2749,N2750,N2751,N2760,N2761,N2766,N2771,N2772,N2773,N2774,
     N2775,N2776,N2777,N2778,N2781,N2782,N2783,N2784,N2789,N2790,
     N2791,N2792,N2793,N2796,N2800,N2803,N2806,N2809,N2810,N2811,
     N2812,N2817,N2820,N2826,N2829,N2830,N2831,N2837,N2838,N2839,
     N2840,N2841,N2844,N2854,N2859,N2869,N2874,N2877,N2880,N2881,
     N2882,N2885,N2888,N2894,N2895,N2896,N2897,N2898,N2899,N2900,
     N2901,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2931,
     N2938,N2939,N2963,N2972,N2975,N2978,N2981,N2984,N2985,N2986,
     N2989,N2992,N2995,N2998,N3001,N3004,N3007,N3008,N3009,N3010,
     N3013,N3016,N3019,N3022,N3025,N3028,N3029,N3030,N3035,N3036,
     N3037,N3039,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3053,
     N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3064,N3065,
     N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,
     N3076,N3088,N3091,N3110,N3113,N3137,N3140,N3143,N3146,N3149,
     N3152,N3157,N3160,N3163,N3166,N3169,N3172,N3175,N3176,N3177,
     N3178,N3180,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,
     N3195,N3196,N3197,N3208,N3215,N3216,N3217,N3218,N3219,N3220,
     N3222,N3223,N3230,N3231,N3238,N3241,N3244,N3247,N3250,N3253,
     N3256,N3259,N3262,N3265,N3268,N3271,N3274,N3277,N3281,N3282,
     N3283,N3284,N3286,N3288,N3289,N3291,N3293,N3295,N3296,N3299,
     N3301,N3302,N3304,N3306,N3308,N3309,N3312,N3314,N3315,N3318,
     N3321,N3324,N3327,N3330,N3333,N3334,N3335,N3336,N3337,N3340,
     N3344,N3348,N3352,N3356,N3360,N3364,N3367,N3370,N3374,N3378,
     N3382,N3386,N3390,N3394,N3397,N3400,N3401,N3402,N3403,N3404,
     N3405,N3406,N3409,N3410,N3412,N3414,N3416,N3418,N3420,N3422,
     N3428,N3430,N3432,N3434,N3436,N3438,N3440,N3450,N3453,N3456,
     N3459,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,
     N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3496,N3498,
     N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,
     N3509,N3510,N3511,N3512,N3513,N3515,N3517,N3522,N3525,N3528,
     N3531,N3534,N3537,N3540,N3543,N3551,N3552,N3553,N3554,N3555,
     N3556,N3557,N3558,N3559,N3563,N3564,N3565,N3566,N3567,N3568,
     N3569,N3570,N3576,N3579,N3585,N3588,N3592,N3593,N3594,N3595,
     N3596,N3597,N3598,N3599,N3600,N3603,N3608,N3612,N3615,N3616,
     N3622,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3640,N3644,
     N3647,N3648,N3654,N3661,N3662,N3667,N3668,N3669,N3670,N3691,
     N3692,N3693,N3694,N3695,N3696,N3697,N3716,N3717,N3718,N3719,
     N3720,N3721,N3722,N3723,N3726,N3727,N3728,N3729,N3730,N3731,
     N3732,N3733,N3734,N3735,N3736,N3737,N3740,N3741,N3742,N3743,
     N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3753,N3754,N3758,
     N3761,N3762,N3767,N3771,N3774,N3775,N3778,N3779,N3780,N3790,
     N3793,N3794,N3802,N3805,N3806,N3807,N3808,N3811,N3812,N3813,
     N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,
     N3826,N3827,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3843,
     N3852,N3857,N3858,N3859,N3864,N3869,N3870,N3876,N3877, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate591inter0, gate591inter1, gate591inter2, gate591inter3, gate591inter4, gate591inter5, gate591inter6, gate591inter7, gate591inter8, gate591inter9, gate591inter10, gate591inter11, gate591inter12, gate1081inter0, gate1081inter1, gate1081inter2, gate1081inter3, gate1081inter4, gate1081inter5, gate1081inter6, gate1081inter7, gate1081inter8, gate1081inter9, gate1081inter10, gate1081inter11, gate1081inter12, gate783inter0, gate783inter1, gate783inter2, gate783inter3, gate783inter4, gate783inter5, gate783inter6, gate783inter7, gate783inter8, gate783inter9, gate783inter10, gate783inter11, gate783inter12, gate1116inter0, gate1116inter1, gate1116inter2, gate1116inter3, gate1116inter4, gate1116inter5, gate1116inter6, gate1116inter7, gate1116inter8, gate1116inter9, gate1116inter10, gate1116inter11, gate1116inter12, gate716inter0, gate716inter1, gate716inter2, gate716inter3, gate716inter4, gate716inter5, gate716inter6, gate716inter7, gate716inter8, gate716inter9, gate716inter10, gate716inter11, gate716inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate651inter0, gate651inter1, gate651inter2, gate651inter3, gate651inter4, gate651inter5, gate651inter6, gate651inter7, gate651inter8, gate651inter9, gate651inter10, gate651inter11, gate651inter12, gate650inter0, gate650inter1, gate650inter2, gate650inter3, gate650inter4, gate650inter5, gate650inter6, gate650inter7, gate650inter8, gate650inter9, gate650inter10, gate650inter11, gate650inter12, gate320inter0, gate320inter1, gate320inter2, gate320inter3, gate320inter4, gate320inter5, gate320inter6, gate320inter7, gate320inter8, gate320inter9, gate320inter10, gate320inter11, gate320inter12, gate587inter0, gate587inter1, gate587inter2, gate587inter3, gate587inter4, gate587inter5, gate587inter6, gate587inter7, gate587inter8, gate587inter9, gate587inter10, gate587inter11, gate587inter12, gate753inter0, gate753inter1, gate753inter2, gate753inter3, gate753inter4, gate753inter5, gate753inter6, gate753inter7, gate753inter8, gate753inter9, gate753inter10, gate753inter11, gate753inter12, gate745inter0, gate745inter1, gate745inter2, gate745inter3, gate745inter4, gate745inter5, gate745inter6, gate745inter7, gate745inter8, gate745inter9, gate745inter10, gate745inter11, gate745inter12, gate532inter0, gate532inter1, gate532inter2, gate532inter3, gate532inter4, gate532inter5, gate532inter6, gate532inter7, gate532inter8, gate532inter9, gate532inter10, gate532inter11, gate532inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate739inter0, gate739inter1, gate739inter2, gate739inter3, gate739inter4, gate739inter5, gate739inter6, gate739inter7, gate739inter8, gate739inter9, gate739inter10, gate739inter11, gate739inter12, gate865inter0, gate865inter1, gate865inter2, gate865inter3, gate865inter4, gate865inter5, gate865inter6, gate865inter7, gate865inter8, gate865inter9, gate865inter10, gate865inter11, gate865inter12, gate300inter0, gate300inter1, gate300inter2, gate300inter3, gate300inter4, gate300inter5, gate300inter6, gate300inter7, gate300inter8, gate300inter9, gate300inter10, gate300inter11, gate300inter12, gate1069inter0, gate1069inter1, gate1069inter2, gate1069inter3, gate1069inter4, gate1069inter5, gate1069inter6, gate1069inter7, gate1069inter8, gate1069inter9, gate1069inter10, gate1069inter11, gate1069inter12, gate555inter0, gate555inter1, gate555inter2, gate555inter3, gate555inter4, gate555inter5, gate555inter6, gate555inter7, gate555inter8, gate555inter9, gate555inter10, gate555inter11, gate555inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate641inter0, gate641inter1, gate641inter2, gate641inter3, gate641inter4, gate641inter5, gate641inter6, gate641inter7, gate641inter8, gate641inter9, gate641inter10, gate641inter11, gate641inter12, gate583inter0, gate583inter1, gate583inter2, gate583inter3, gate583inter4, gate583inter5, gate583inter6, gate583inter7, gate583inter8, gate583inter9, gate583inter10, gate583inter11, gate583inter12, gate1079inter0, gate1079inter1, gate1079inter2, gate1079inter3, gate1079inter4, gate1079inter5, gate1079inter6, gate1079inter7, gate1079inter8, gate1079inter9, gate1079inter10, gate1079inter11, gate1079inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate1141inter0, gate1141inter1, gate1141inter2, gate1141inter3, gate1141inter4, gate1141inter5, gate1141inter6, gate1141inter7, gate1141inter8, gate1141inter9, gate1141inter10, gate1141inter11, gate1141inter12, gate538inter0, gate538inter1, gate538inter2, gate538inter3, gate538inter4, gate538inter5, gate538inter6, gate538inter7, gate538inter8, gate538inter9, gate538inter10, gate538inter11, gate538inter12, gate646inter0, gate646inter1, gate646inter2, gate646inter3, gate646inter4, gate646inter5, gate646inter6, gate646inter7, gate646inter8, gate646inter9, gate646inter10, gate646inter11, gate646inter12, gate1051inter0, gate1051inter1, gate1051inter2, gate1051inter3, gate1051inter4, gate1051inter5, gate1051inter6, gate1051inter7, gate1051inter8, gate1051inter9, gate1051inter10, gate1051inter11, gate1051inter12, gate1105inter0, gate1105inter1, gate1105inter2, gate1105inter3, gate1105inter4, gate1105inter5, gate1105inter6, gate1105inter7, gate1105inter8, gate1105inter9, gate1105inter10, gate1105inter11, gate1105inter12, gate1056inter0, gate1056inter1, gate1056inter2, gate1056inter3, gate1056inter4, gate1056inter5, gate1056inter6, gate1056inter7, gate1056inter8, gate1056inter9, gate1056inter10, gate1056inter11, gate1056inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate647inter0, gate647inter1, gate647inter2, gate647inter3, gate647inter4, gate647inter5, gate647inter6, gate647inter7, gate647inter8, gate647inter9, gate647inter10, gate647inter11, gate647inter12, gate1182inter0, gate1182inter1, gate1182inter2, gate1182inter3, gate1182inter4, gate1182inter5, gate1182inter6, gate1182inter7, gate1182inter8, gate1182inter9, gate1182inter10, gate1182inter11, gate1182inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate930inter0, gate930inter1, gate930inter2, gate930inter3, gate930inter4, gate930inter5, gate930inter6, gate930inter7, gate930inter8, gate930inter9, gate930inter10, gate930inter11, gate930inter12, gate1126inter0, gate1126inter1, gate1126inter2, gate1126inter3, gate1126inter4, gate1126inter5, gate1126inter6, gate1126inter7, gate1126inter8, gate1126inter9, gate1126inter10, gate1126inter11, gate1126inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate736inter0, gate736inter1, gate736inter2, gate736inter3, gate736inter4, gate736inter5, gate736inter6, gate736inter7, gate736inter8, gate736inter9, gate736inter10, gate736inter11, gate736inter12, gate638inter0, gate638inter1, gate638inter2, gate638inter3, gate638inter4, gate638inter5, gate638inter6, gate638inter7, gate638inter8, gate638inter9, gate638inter10, gate638inter11, gate638inter12, gate1169inter0, gate1169inter1, gate1169inter2, gate1169inter3, gate1169inter4, gate1169inter5, gate1169inter6, gate1169inter7, gate1169inter8, gate1169inter9, gate1169inter10, gate1169inter11, gate1169inter12, gate644inter0, gate644inter1, gate644inter2, gate644inter3, gate644inter4, gate644inter5, gate644inter6, gate644inter7, gate644inter8, gate644inter9, gate644inter10, gate644inter11, gate644inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate883inter0, gate883inter1, gate883inter2, gate883inter3, gate883inter4, gate883inter5, gate883inter6, gate883inter7, gate883inter8, gate883inter9, gate883inter10, gate883inter11, gate883inter12, gate536inter0, gate536inter1, gate536inter2, gate536inter3, gate536inter4, gate536inter5, gate536inter6, gate536inter7, gate536inter8, gate536inter9, gate536inter10, gate536inter11, gate536inter12, gate534inter0, gate534inter1, gate534inter2, gate534inter3, gate534inter4, gate534inter5, gate534inter6, gate534inter7, gate534inter8, gate534inter9, gate534inter10, gate534inter11, gate534inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate609inter0, gate609inter1, gate609inter2, gate609inter3, gate609inter4, gate609inter5, gate609inter6, gate609inter7, gate609inter8, gate609inter9, gate609inter10, gate609inter11, gate609inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate884inter0, gate884inter1, gate884inter2, gate884inter3, gate884inter4, gate884inter5, gate884inter6, gate884inter7, gate884inter8, gate884inter9, gate884inter10, gate884inter11, gate884inter12, gate558inter0, gate558inter1, gate558inter2, gate558inter3, gate558inter4, gate558inter5, gate558inter6, gate558inter7, gate558inter8, gate558inter9, gate558inter10, gate558inter11, gate558inter12, gate586inter0, gate586inter1, gate586inter2, gate586inter3, gate586inter4, gate586inter5, gate586inter6, gate586inter7, gate586inter8, gate586inter9, gate586inter10, gate586inter11, gate586inter12, gate885inter0, gate885inter1, gate885inter2, gate885inter3, gate885inter4, gate885inter5, gate885inter6, gate885inter7, gate885inter8, gate885inter9, gate885inter10, gate885inter11, gate885inter12, gate777inter0, gate777inter1, gate777inter2, gate777inter3, gate777inter4, gate777inter5, gate777inter6, gate777inter7, gate777inter8, gate777inter9, gate777inter10, gate777inter11, gate777inter12;



buf1 gate1( .a(N219), .O(N398) );
buf1 gate2( .a(N219), .O(N400) );
buf1 gate3( .a(N219), .O(N401) );
and2 gate4( .a(N1), .b(N3), .O(N405) );
inv1 gate5( .a(N230), .O(N408) );
buf1 gate6( .a(N253), .O(N419) );
buf1 gate7( .a(N253), .O(N420) );
inv1 gate8( .a(N262), .O(N425) );
buf1 gate9( .a(N290), .O(N456) );
buf1 gate10( .a(N290), .O(N457) );
buf1 gate11( .a(N290), .O(N458) );
and4 gate12( .a(N309), .b(N305), .c(N301), .d(N297), .O(N485) );
inv1 gate13( .a(N405), .O(N486) );
inv1 gate14( .a(N44), .O(N487) );
inv1 gate15( .a(N132), .O(N488) );
inv1 gate16( .a(N82), .O(N489) );
inv1 gate17( .a(N96), .O(N490) );
inv1 gate18( .a(N69), .O(N491) );
inv1 gate19( .a(N120), .O(N492) );
inv1 gate20( .a(N57), .O(N493) );
inv1 gate21( .a(N108), .O(N494) );
and3 gate22( .a(N2), .b(N15), .c(N237), .O(N495) );
buf1 gate23( .a(N237), .O(N496) );
and2 gate24( .a(N37), .b(N37), .O(N499) );
buf1 gate25( .a(N219), .O(N500) );
buf1 gate26( .a(N8), .O(N503) );
buf1 gate27( .a(N8), .O(N506) );
buf1 gate28( .a(N227), .O(N509) );
buf1 gate29( .a(N234), .O(N521) );
inv1 gate30( .a(N241), .O(N533) );
inv1 gate31( .a(N246), .O(N537) );
and2 gate32( .a(N11), .b(N246), .O(N543) );
and4 gate33( .a(N132), .b(N82), .c(N96), .d(N44), .O(N544) );
and4 gate34( .a(N120), .b(N57), .c(N108), .d(N69), .O(N547) );
buf1 gate35( .a(N227), .O(N550) );
buf1 gate36( .a(N234), .O(N562) );
inv1 gate37( .a(N256), .O(N574) );
inv1 gate38( .a(N259), .O(N578) );
buf1 gate39( .a(N319), .O(N582) );
buf1 gate40( .a(N322), .O(N594) );
inv1 gate41( .a(N328), .O(N606) );
inv1 gate42( .a(N331), .O(N607) );
inv1 gate43( .a(N334), .O(N608) );
inv1 gate44( .a(N337), .O(N609) );
inv1 gate45( .a(N340), .O(N610) );
inv1 gate46( .a(N343), .O(N611) );
inv1 gate47( .a(N352), .O(N612) );
buf1 gate48( .a(N319), .O(N613) );
buf1 gate49( .a(N322), .O(N625) );
buf1 gate50( .a(N16), .O(N637) );
buf1 gate51( .a(N16), .O(N643) );
inv1 gate52( .a(N355), .O(N650) );
and2 gate53( .a(N7), .b(N237), .O(N651) );
inv1 gate54( .a(N263), .O(N655) );
inv1 gate55( .a(N266), .O(N659) );
inv1 gate56( .a(N269), .O(N663) );
inv1 gate57( .a(N272), .O(N667) );
inv1 gate58( .a(N275), .O(N671) );
inv1 gate59( .a(N278), .O(N675) );
inv1 gate60( .a(N281), .O(N679) );
inv1 gate61( .a(N284), .O(N683) );
inv1 gate62( .a(N287), .O(N687) );
buf1 gate63( .a(N29), .O(N693) );
buf1 gate64( .a(N29), .O(N699) );
inv1 gate65( .a(N294), .O(N705) );
inv1 gate66( .a(N297), .O(N711) );
inv1 gate67( .a(N301), .O(N715) );
inv1 gate68( .a(N305), .O(N719) );
inv1 gate69( .a(N309), .O(N723) );
inv1 gate70( .a(N313), .O(N727) );
inv1 gate71( .a(N316), .O(N730) );
inv1 gate72( .a(N346), .O(N733) );
inv1 gate73( .a(N349), .O(N734) );
buf1 gate74( .a(N259), .O(N735) );
buf1 gate75( .a(N256), .O(N738) );
buf1 gate76( .a(N263), .O(N741) );
buf1 gate77( .a(N269), .O(N744) );
buf1 gate78( .a(N266), .O(N747) );
buf1 gate79( .a(N275), .O(N750) );
buf1 gate80( .a(N272), .O(N753) );
buf1 gate81( .a(N281), .O(N756) );
buf1 gate82( .a(N278), .O(N759) );
buf1 gate83( .a(N287), .O(N762) );
buf1 gate84( .a(N284), .O(N765) );
buf1 gate85( .a(N294), .O(N768) );
buf1 gate86( .a(N301), .O(N771) );
buf1 gate87( .a(N297), .O(N774) );
buf1 gate88( .a(N309), .O(N777) );
buf1 gate89( .a(N305), .O(N780) );
buf1 gate90( .a(N316), .O(N783) );
buf1 gate91( .a(N313), .O(N786) );
inv1 gate92( .a(N485), .O(N792) );
inv1 gate93( .a(N495), .O(N799) );
inv1 gate94( .a(N499), .O(N800) );
buf1 gate95( .a(N500), .O(N805) );
nand2 gate96( .a(N331), .b(N606), .O(N900) );
nand2 gate97( .a(N328), .b(N607), .O(N901) );
nand2 gate98( .a(N337), .b(N608), .O(N902) );
nand2 gate99( .a(N334), .b(N609), .O(N903) );

  xor2  gate1620(.a(N610), .b(N343), .O(gate100inter0));
  nand2 gate1621(.a(gate100inter0), .b(s_50), .O(gate100inter1));
  and2  gate1622(.a(N610), .b(N343), .O(gate100inter2));
  inv1  gate1623(.a(s_50), .O(gate100inter3));
  inv1  gate1624(.a(s_51), .O(gate100inter4));
  nand2 gate1625(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1626(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1627(.a(N343), .O(gate100inter7));
  inv1  gate1628(.a(N610), .O(gate100inter8));
  nand2 gate1629(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1630(.a(s_51), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1631(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1632(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1633(.a(gate100inter12), .b(gate100inter1), .O(N904));

  xor2  gate1970(.a(N611), .b(N340), .O(gate101inter0));
  nand2 gate1971(.a(gate101inter0), .b(s_100), .O(gate101inter1));
  and2  gate1972(.a(N611), .b(N340), .O(gate101inter2));
  inv1  gate1973(.a(s_100), .O(gate101inter3));
  inv1  gate1974(.a(s_101), .O(gate101inter4));
  nand2 gate1975(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1976(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1977(.a(N340), .O(gate101inter7));
  inv1  gate1978(.a(N611), .O(gate101inter8));
  nand2 gate1979(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1980(.a(s_101), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1981(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1982(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1983(.a(gate101inter12), .b(gate101inter1), .O(N905));
nand2 gate102( .a(N349), .b(N733), .O(N998) );

  xor2  gate1284(.a(N734), .b(N346), .O(gate103inter0));
  nand2 gate1285(.a(gate103inter0), .b(s_2), .O(gate103inter1));
  and2  gate1286(.a(N734), .b(N346), .O(gate103inter2));
  inv1  gate1287(.a(s_2), .O(gate103inter3));
  inv1  gate1288(.a(s_3), .O(gate103inter4));
  nand2 gate1289(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1290(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1291(.a(N346), .O(gate103inter7));
  inv1  gate1292(.a(N734), .O(gate103inter8));
  nand2 gate1293(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1294(.a(s_3), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1295(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1296(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1297(.a(gate103inter12), .b(gate103inter1), .O(N999));
and2 gate104( .a(N94), .b(N500), .O(N1026) );
and2 gate105( .a(N325), .b(N651), .O(N1027) );
inv1 gate106( .a(N651), .O(N1028) );
nand2 gate107( .a(N231), .b(N651), .O(N1029) );
inv1 gate108( .a(N544), .O(N1032) );
inv1 gate109( .a(N547), .O(N1033) );
and2 gate110( .a(N547), .b(N544), .O(N1034) );
buf1 gate111( .a(N503), .O(N1037) );
inv1 gate112( .a(N509), .O(N1042) );
inv1 gate113( .a(N521), .O(N1053) );
and3 gate114( .a(N80), .b(N509), .c(N521), .O(N1064) );
and3 gate115( .a(N68), .b(N509), .c(N521), .O(N1065) );
and3 gate116( .a(N79), .b(N509), .c(N521), .O(N1066) );
and3 gate117( .a(N78), .b(N509), .c(N521), .O(N1067) );
and3 gate118( .a(N77), .b(N509), .c(N521), .O(N1068) );
and2 gate119( .a(N11), .b(N537), .O(N1069) );
buf1 gate120( .a(N503), .O(N1070) );
inv1 gate121( .a(N550), .O(N1075) );
inv1 gate122( .a(N562), .O(N1086) );
and3 gate123( .a(N76), .b(N550), .c(N562), .O(N1097) );
and3 gate124( .a(N75), .b(N550), .c(N562), .O(N1098) );
and3 gate125( .a(N74), .b(N550), .c(N562), .O(N1099) );
and3 gate126( .a(N73), .b(N550), .c(N562), .O(N1100) );
and3 gate127( .a(N72), .b(N550), .c(N562), .O(N1101) );
inv1 gate128( .a(N582), .O(N1102) );
inv1 gate129( .a(N594), .O(N1113) );
and3 gate130( .a(N114), .b(N582), .c(N594), .O(N1124) );
and3 gate131( .a(N113), .b(N582), .c(N594), .O(N1125) );
and3 gate132( .a(N112), .b(N582), .c(N594), .O(N1126) );
and3 gate133( .a(N111), .b(N582), .c(N594), .O(N1127) );
and2 gate134( .a(N582), .b(N594), .O(N1128) );
nand2 gate135( .a(N900), .b(N901), .O(N1129) );

  xor2  gate1480(.a(N903), .b(N902), .O(gate136inter0));
  nand2 gate1481(.a(gate136inter0), .b(s_30), .O(gate136inter1));
  and2  gate1482(.a(N903), .b(N902), .O(gate136inter2));
  inv1  gate1483(.a(s_30), .O(gate136inter3));
  inv1  gate1484(.a(s_31), .O(gate136inter4));
  nand2 gate1485(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1486(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1487(.a(N902), .O(gate136inter7));
  inv1  gate1488(.a(N903), .O(gate136inter8));
  nand2 gate1489(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1490(.a(s_31), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1491(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1492(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1493(.a(gate136inter12), .b(gate136inter1), .O(N1133));
nand2 gate137( .a(N904), .b(N905), .O(N1137) );
inv1 gate138( .a(N741), .O(N1140) );

  xor2  gate1368(.a(N612), .b(N741), .O(gate139inter0));
  nand2 gate1369(.a(gate139inter0), .b(s_14), .O(gate139inter1));
  and2  gate1370(.a(N612), .b(N741), .O(gate139inter2));
  inv1  gate1371(.a(s_14), .O(gate139inter3));
  inv1  gate1372(.a(s_15), .O(gate139inter4));
  nand2 gate1373(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1374(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1375(.a(N741), .O(gate139inter7));
  inv1  gate1376(.a(N612), .O(gate139inter8));
  nand2 gate1377(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1378(.a(s_15), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1379(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1380(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1381(.a(gate139inter12), .b(gate139inter1), .O(N1141));
inv1 gate140( .a(N744), .O(N1142) );
inv1 gate141( .a(N747), .O(N1143) );
inv1 gate142( .a(N750), .O(N1144) );
inv1 gate143( .a(N753), .O(N1145) );
inv1 gate144( .a(N613), .O(N1146) );
inv1 gate145( .a(N625), .O(N1157) );
and3 gate146( .a(N118), .b(N613), .c(N625), .O(N1168) );
and3 gate147( .a(N107), .b(N613), .c(N625), .O(N1169) );
and3 gate148( .a(N117), .b(N613), .c(N625), .O(N1170) );
and3 gate149( .a(N116), .b(N613), .c(N625), .O(N1171) );
and3 gate150( .a(N115), .b(N613), .c(N625), .O(N1172) );
inv1 gate151( .a(N637), .O(N1173) );
inv1 gate152( .a(N643), .O(N1178) );
inv1 gate153( .a(N768), .O(N1184) );
nand2 gate154( .a(N768), .b(N650), .O(N1185) );
inv1 gate155( .a(N771), .O(N1186) );
inv1 gate156( .a(N774), .O(N1187) );
inv1 gate157( .a(N777), .O(N1188) );
inv1 gate158( .a(N780), .O(N1189) );
buf1 gate159( .a(N506), .O(N1190) );
buf1 gate160( .a(N506), .O(N1195) );
inv1 gate161( .a(N693), .O(N1200) );
inv1 gate162( .a(N699), .O(N1205) );
inv1 gate163( .a(N735), .O(N1210) );
inv1 gate164( .a(N738), .O(N1211) );
inv1 gate165( .a(N756), .O(N1212) );
inv1 gate166( .a(N759), .O(N1213) );
inv1 gate167( .a(N762), .O(N1214) );
inv1 gate168( .a(N765), .O(N1215) );
nand2 gate169( .a(N998), .b(N999), .O(N1216) );
buf1 gate170( .a(N574), .O(N1219) );
buf1 gate171( .a(N578), .O(N1222) );
buf1 gate172( .a(N655), .O(N1225) );
buf1 gate173( .a(N659), .O(N1228) );
buf1 gate174( .a(N663), .O(N1231) );
buf1 gate175( .a(N667), .O(N1234) );
buf1 gate176( .a(N671), .O(N1237) );
buf1 gate177( .a(N675), .O(N1240) );
buf1 gate178( .a(N679), .O(N1243) );
buf1 gate179( .a(N683), .O(N1246) );
inv1 gate180( .a(N783), .O(N1249) );
inv1 gate181( .a(N786), .O(N1250) );
buf1 gate182( .a(N687), .O(N1251) );
buf1 gate183( .a(N705), .O(N1254) );
buf1 gate184( .a(N711), .O(N1257) );
buf1 gate185( .a(N715), .O(N1260) );
buf1 gate186( .a(N719), .O(N1263) );
buf1 gate187( .a(N723), .O(N1266) );
inv1 gate188( .a(N1027), .O(N1269) );
and2 gate189( .a(N325), .b(N1032), .O(N1275) );
and2 gate190( .a(N231), .b(N1033), .O(N1276) );
buf1 gate191( .a(N1034), .O(N1277) );
or2 gate192( .a(N1069), .b(N543), .O(N1302) );
nand2 gate193( .a(N352), .b(N1140), .O(N1351) );
nand2 gate194( .a(N747), .b(N1142), .O(N1352) );
nand2 gate195( .a(N744), .b(N1143), .O(N1353) );
nand2 gate196( .a(N753), .b(N1144), .O(N1354) );
nand2 gate197( .a(N750), .b(N1145), .O(N1355) );
nand2 gate198( .a(N355), .b(N1184), .O(N1395) );

  xor2  gate1270(.a(N1186), .b(N774), .O(gate199inter0));
  nand2 gate1271(.a(gate199inter0), .b(s_0), .O(gate199inter1));
  and2  gate1272(.a(N1186), .b(N774), .O(gate199inter2));
  inv1  gate1273(.a(s_0), .O(gate199inter3));
  inv1  gate1274(.a(s_1), .O(gate199inter4));
  nand2 gate1275(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1276(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1277(.a(N774), .O(gate199inter7));
  inv1  gate1278(.a(N1186), .O(gate199inter8));
  nand2 gate1279(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1280(.a(s_1), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1281(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1282(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1283(.a(gate199inter12), .b(gate199inter1), .O(N1396));
nand2 gate200( .a(N771), .b(N1187), .O(N1397) );
nand2 gate201( .a(N780), .b(N1188), .O(N1398) );
nand2 gate202( .a(N777), .b(N1189), .O(N1399) );
nand2 gate203( .a(N738), .b(N1210), .O(N1422) );
nand2 gate204( .a(N735), .b(N1211), .O(N1423) );
nand2 gate205( .a(N759), .b(N1212), .O(N1424) );

  xor2  gate1802(.a(N1213), .b(N756), .O(gate206inter0));
  nand2 gate1803(.a(gate206inter0), .b(s_76), .O(gate206inter1));
  and2  gate1804(.a(N1213), .b(N756), .O(gate206inter2));
  inv1  gate1805(.a(s_76), .O(gate206inter3));
  inv1  gate1806(.a(s_77), .O(gate206inter4));
  nand2 gate1807(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1808(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1809(.a(N756), .O(gate206inter7));
  inv1  gate1810(.a(N1213), .O(gate206inter8));
  nand2 gate1811(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1812(.a(s_77), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1813(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1814(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1815(.a(gate206inter12), .b(gate206inter1), .O(N1425));
nand2 gate207( .a(N765), .b(N1214), .O(N1426) );

  xor2  gate1942(.a(N1215), .b(N762), .O(gate208inter0));
  nand2 gate1943(.a(gate208inter0), .b(s_96), .O(gate208inter1));
  and2  gate1944(.a(N1215), .b(N762), .O(gate208inter2));
  inv1  gate1945(.a(s_96), .O(gate208inter3));
  inv1  gate1946(.a(s_97), .O(gate208inter4));
  nand2 gate1947(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1948(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1949(.a(N762), .O(gate208inter7));
  inv1  gate1950(.a(N1215), .O(gate208inter8));
  nand2 gate1951(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1952(.a(s_97), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1953(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1954(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1955(.a(gate208inter12), .b(gate208inter1), .O(N1427));
nand2 gate209( .a(N786), .b(N1249), .O(N1440) );

  xor2  gate1886(.a(N1250), .b(N783), .O(gate210inter0));
  nand2 gate1887(.a(gate210inter0), .b(s_88), .O(gate210inter1));
  and2  gate1888(.a(N1250), .b(N783), .O(gate210inter2));
  inv1  gate1889(.a(s_88), .O(gate210inter3));
  inv1  gate1890(.a(s_89), .O(gate210inter4));
  nand2 gate1891(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1892(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1893(.a(N783), .O(gate210inter7));
  inv1  gate1894(.a(N1250), .O(gate210inter8));
  nand2 gate1895(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1896(.a(s_89), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1897(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1898(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1899(.a(gate210inter12), .b(gate210inter1), .O(N1441));
inv1 gate211( .a(N1034), .O(N1448) );
inv1 gate212( .a(N1275), .O(N1449) );
inv1 gate213( .a(N1276), .O(N1450) );
and3 gate214( .a(N93), .b(N1042), .c(N1053), .O(N1451) );
and3 gate215( .a(N55), .b(N509), .c(N1053), .O(N1452) );
and3 gate216( .a(N67), .b(N1042), .c(N521), .O(N1453) );
and3 gate217( .a(N81), .b(N1042), .c(N1053), .O(N1454) );
and3 gate218( .a(N43), .b(N509), .c(N1053), .O(N1455) );
and3 gate219( .a(N56), .b(N1042), .c(N521), .O(N1456) );
and3 gate220( .a(N92), .b(N1042), .c(N1053), .O(N1457) );
and3 gate221( .a(N54), .b(N509), .c(N1053), .O(N1458) );
and3 gate222( .a(N66), .b(N1042), .c(N521), .O(N1459) );
and3 gate223( .a(N91), .b(N1042), .c(N1053), .O(N1460) );
and3 gate224( .a(N53), .b(N509), .c(N1053), .O(N1461) );
and3 gate225( .a(N65), .b(N1042), .c(N521), .O(N1462) );
and3 gate226( .a(N90), .b(N1042), .c(N1053), .O(N1463) );
and3 gate227( .a(N52), .b(N509), .c(N1053), .O(N1464) );
and3 gate228( .a(N64), .b(N1042), .c(N521), .O(N1465) );
and3 gate229( .a(N89), .b(N1075), .c(N1086), .O(N1466) );
and3 gate230( .a(N51), .b(N550), .c(N1086), .O(N1467) );
and3 gate231( .a(N63), .b(N1075), .c(N562), .O(N1468) );
and3 gate232( .a(N88), .b(N1075), .c(N1086), .O(N1469) );
and3 gate233( .a(N50), .b(N550), .c(N1086), .O(N1470) );
and3 gate234( .a(N62), .b(N1075), .c(N562), .O(N1471) );
and3 gate235( .a(N87), .b(N1075), .c(N1086), .O(N1472) );
and3 gate236( .a(N49), .b(N550), .c(N1086), .O(N1473) );
and2 gate237( .a(N1075), .b(N562), .O(N1474) );
and3 gate238( .a(N86), .b(N1075), .c(N1086), .O(N1475) );
and3 gate239( .a(N48), .b(N550), .c(N1086), .O(N1476) );
and3 gate240( .a(N61), .b(N1075), .c(N562), .O(N1477) );
and3 gate241( .a(N85), .b(N1075), .c(N1086), .O(N1478) );
and3 gate242( .a(N47), .b(N550), .c(N1086), .O(N1479) );
and3 gate243( .a(N60), .b(N1075), .c(N562), .O(N1480) );
and3 gate244( .a(N138), .b(N1102), .c(N1113), .O(N1481) );
and3 gate245( .a(N102), .b(N582), .c(N1113), .O(N1482) );
and3 gate246( .a(N126), .b(N1102), .c(N594), .O(N1483) );
and3 gate247( .a(N137), .b(N1102), .c(N1113), .O(N1484) );
and3 gate248( .a(N101), .b(N582), .c(N1113), .O(N1485) );
and3 gate249( .a(N125), .b(N1102), .c(N594), .O(N1486) );
and3 gate250( .a(N136), .b(N1102), .c(N1113), .O(N1487) );
and3 gate251( .a(N100), .b(N582), .c(N1113), .O(N1488) );
and3 gate252( .a(N124), .b(N1102), .c(N594), .O(N1489) );
and3 gate253( .a(N135), .b(N1102), .c(N1113), .O(N1490) );
and3 gate254( .a(N99), .b(N582), .c(N1113), .O(N1491) );
and3 gate255( .a(N123), .b(N1102), .c(N594), .O(N1492) );
and2 gate256( .a(N1102), .b(N1113), .O(N1493) );
and2 gate257( .a(N582), .b(N1113), .O(N1494) );
and2 gate258( .a(N1102), .b(N594), .O(N1495) );
inv1 gate259( .a(N1129), .O(N1496) );
inv1 gate260( .a(N1133), .O(N1499) );
nand2 gate261( .a(N1351), .b(N1141), .O(N1502) );
nand2 gate262( .a(N1352), .b(N1353), .O(N1506) );
nand2 gate263( .a(N1354), .b(N1355), .O(N1510) );
buf1 gate264( .a(N1137), .O(N1513) );
buf1 gate265( .a(N1137), .O(N1516) );
inv1 gate266( .a(N1219), .O(N1519) );
inv1 gate267( .a(N1222), .O(N1520) );
inv1 gate268( .a(N1225), .O(N1521) );
inv1 gate269( .a(N1228), .O(N1522) );
inv1 gate270( .a(N1231), .O(N1523) );
inv1 gate271( .a(N1234), .O(N1524) );
inv1 gate272( .a(N1237), .O(N1525) );
inv1 gate273( .a(N1240), .O(N1526) );
inv1 gate274( .a(N1243), .O(N1527) );
inv1 gate275( .a(N1246), .O(N1528) );
and3 gate276( .a(N142), .b(N1146), .c(N1157), .O(N1529) );
and3 gate277( .a(N106), .b(N613), .c(N1157), .O(N1530) );
and3 gate278( .a(N130), .b(N1146), .c(N625), .O(N1531) );
and3 gate279( .a(N131), .b(N1146), .c(N1157), .O(N1532) );
and3 gate280( .a(N95), .b(N613), .c(N1157), .O(N1533) );
and3 gate281( .a(N119), .b(N1146), .c(N625), .O(N1534) );
and3 gate282( .a(N141), .b(N1146), .c(N1157), .O(N1535) );
and3 gate283( .a(N105), .b(N613), .c(N1157), .O(N1536) );
and3 gate284( .a(N129), .b(N1146), .c(N625), .O(N1537) );
and3 gate285( .a(N140), .b(N1146), .c(N1157), .O(N1538) );
and3 gate286( .a(N104), .b(N613), .c(N1157), .O(N1539) );
and3 gate287( .a(N128), .b(N1146), .c(N625), .O(N1540) );
and3 gate288( .a(N139), .b(N1146), .c(N1157), .O(N1541) );
and3 gate289( .a(N103), .b(N613), .c(N1157), .O(N1542) );
and3 gate290( .a(N127), .b(N1146), .c(N625), .O(N1543) );
and2 gate291( .a(N19), .b(N1173), .O(N1544) );
and2 gate292( .a(N4), .b(N1173), .O(N1545) );
and2 gate293( .a(N20), .b(N1173), .O(N1546) );
and2 gate294( .a(N5), .b(N1173), .O(N1547) );
and2 gate295( .a(N21), .b(N1178), .O(N1548) );
and2 gate296( .a(N22), .b(N1178), .O(N1549) );
and2 gate297( .a(N23), .b(N1178), .O(N1550) );
and2 gate298( .a(N6), .b(N1178), .O(N1551) );
and2 gate299( .a(N24), .b(N1178), .O(N1552) );

  xor2  gate1522(.a(N1185), .b(N1395), .O(gate300inter0));
  nand2 gate1523(.a(gate300inter0), .b(s_36), .O(gate300inter1));
  and2  gate1524(.a(N1185), .b(N1395), .O(gate300inter2));
  inv1  gate1525(.a(s_36), .O(gate300inter3));
  inv1  gate1526(.a(s_37), .O(gate300inter4));
  nand2 gate1527(.a(gate300inter4), .b(gate300inter3), .O(gate300inter5));
  nor2  gate1528(.a(gate300inter5), .b(gate300inter2), .O(gate300inter6));
  inv1  gate1529(.a(N1395), .O(gate300inter7));
  inv1  gate1530(.a(N1185), .O(gate300inter8));
  nand2 gate1531(.a(gate300inter8), .b(gate300inter7), .O(gate300inter9));
  nand2 gate1532(.a(s_37), .b(gate300inter3), .O(gate300inter10));
  nor2  gate1533(.a(gate300inter10), .b(gate300inter9), .O(gate300inter11));
  nor2  gate1534(.a(gate300inter11), .b(gate300inter6), .O(gate300inter12));
  nand2 gate1535(.a(gate300inter12), .b(gate300inter1), .O(N1553));
nand2 gate301( .a(N1396), .b(N1397), .O(N1557) );
nand2 gate302( .a(N1398), .b(N1399), .O(N1561) );
and2 gate303( .a(N25), .b(N1200), .O(N1564) );
and2 gate304( .a(N32), .b(N1200), .O(N1565) );
and2 gate305( .a(N26), .b(N1200), .O(N1566) );
and2 gate306( .a(N33), .b(N1200), .O(N1567) );
and2 gate307( .a(N27), .b(N1205), .O(N1568) );
and2 gate308( .a(N34), .b(N1205), .O(N1569) );
and2 gate309( .a(N35), .b(N1205), .O(N1570) );
and2 gate310( .a(N28), .b(N1205), .O(N1571) );
inv1 gate311( .a(N1251), .O(N1572) );
inv1 gate312( .a(N1254), .O(N1573) );
inv1 gate313( .a(N1257), .O(N1574) );
inv1 gate314( .a(N1260), .O(N1575) );
inv1 gate315( .a(N1263), .O(N1576) );
inv1 gate316( .a(N1266), .O(N1577) );
nand2 gate317( .a(N1422), .b(N1423), .O(N1578) );
inv1 gate318( .a(N1216), .O(N1581) );
nand2 gate319( .a(N1426), .b(N1427), .O(N1582) );

  xor2  gate1410(.a(N1425), .b(N1424), .O(gate320inter0));
  nand2 gate1411(.a(gate320inter0), .b(s_20), .O(gate320inter1));
  and2  gate1412(.a(N1425), .b(N1424), .O(gate320inter2));
  inv1  gate1413(.a(s_20), .O(gate320inter3));
  inv1  gate1414(.a(s_21), .O(gate320inter4));
  nand2 gate1415(.a(gate320inter4), .b(gate320inter3), .O(gate320inter5));
  nor2  gate1416(.a(gate320inter5), .b(gate320inter2), .O(gate320inter6));
  inv1  gate1417(.a(N1424), .O(gate320inter7));
  inv1  gate1418(.a(N1425), .O(gate320inter8));
  nand2 gate1419(.a(gate320inter8), .b(gate320inter7), .O(gate320inter9));
  nand2 gate1420(.a(s_21), .b(gate320inter3), .O(gate320inter10));
  nor2  gate1421(.a(gate320inter10), .b(gate320inter9), .O(gate320inter11));
  nor2  gate1422(.a(gate320inter11), .b(gate320inter6), .O(gate320inter12));
  nand2 gate1423(.a(gate320inter12), .b(gate320inter1), .O(N1585));
nand2 gate321( .a(N1440), .b(N1441), .O(N1588) );
and2 gate322( .a(N1449), .b(N1450), .O(N1591) );
or4 gate323( .a(N1451), .b(N1452), .c(N1453), .d(N1064), .O(N1596) );
or4 gate324( .a(N1454), .b(N1455), .c(N1456), .d(N1065), .O(N1600) );
or4 gate325( .a(N1457), .b(N1458), .c(N1459), .d(N1066), .O(N1606) );
or4 gate326( .a(N1460), .b(N1461), .c(N1462), .d(N1067), .O(N1612) );
or4 gate327( .a(N1463), .b(N1464), .c(N1465), .d(N1068), .O(N1615) );
or4 gate328( .a(N1466), .b(N1467), .c(N1468), .d(N1097), .O(N1619) );
or4 gate329( .a(N1469), .b(N1470), .c(N1471), .d(N1098), .O(N1624) );
or4 gate330( .a(N1472), .b(N1473), .c(N1474), .d(N1099), .O(N1628) );
or4 gate331( .a(N1475), .b(N1476), .c(N1477), .d(N1100), .O(N1631) );
or4 gate332( .a(N1478), .b(N1479), .c(N1480), .d(N1101), .O(N1634) );
or4 gate333( .a(N1481), .b(N1482), .c(N1483), .d(N1124), .O(N1637) );
or4 gate334( .a(N1484), .b(N1485), .c(N1486), .d(N1125), .O(N1642) );
or4 gate335( .a(N1487), .b(N1488), .c(N1489), .d(N1126), .O(N1647) );
or4 gate336( .a(N1490), .b(N1491), .c(N1492), .d(N1127), .O(N1651) );
or4 gate337( .a(N1493), .b(N1494), .c(N1495), .d(N1128), .O(N1656) );
or4 gate338( .a(N1532), .b(N1533), .c(N1534), .d(N1169), .O(N1676) );
or4 gate339( .a(N1535), .b(N1536), .c(N1537), .d(N1170), .O(N1681) );
or4 gate340( .a(N1538), .b(N1539), .c(N1540), .d(N1171), .O(N1686) );
or4 gate341( .a(N1541), .b(N1542), .c(N1543), .d(N1172), .O(N1690) );
or4 gate342( .a(N1529), .b(N1530), .c(N1531), .d(N1168), .O(N1708) );
buf1 gate343( .a(N1591), .O(N1726) );
inv1 gate344( .a(N1502), .O(N1770) );
inv1 gate345( .a(N1506), .O(N1773) );
inv1 gate346( .a(N1513), .O(N1776) );
inv1 gate347( .a(N1516), .O(N1777) );
buf1 gate348( .a(N1510), .O(N1778) );
buf1 gate349( .a(N1510), .O(N1781) );
and3 gate350( .a(N1133), .b(N1129), .c(N1513), .O(N1784) );
and3 gate351( .a(N1499), .b(N1496), .c(N1516), .O(N1785) );
inv1 gate352( .a(N1553), .O(N1795) );
inv1 gate353( .a(N1557), .O(N1798) );
buf1 gate354( .a(N1561), .O(N1801) );
buf1 gate355( .a(N1561), .O(N1804) );
inv1 gate356( .a(N1588), .O(N1807) );
inv1 gate357( .a(N1578), .O(N1808) );
nand2 gate358( .a(N1578), .b(N1581), .O(N1809) );
inv1 gate359( .a(N1582), .O(N1810) );
inv1 gate360( .a(N1585), .O(N1811) );
and2 gate361( .a(N1596), .b(N241), .O(N1813) );
and2 gate362( .a(N1606), .b(N241), .O(N1814) );
and2 gate363( .a(N1600), .b(N241), .O(N1815) );
inv1 gate364( .a(N1642), .O(N1816) );
inv1 gate365( .a(N1647), .O(N1817) );
inv1 gate366( .a(N1637), .O(N1818) );
inv1 gate367( .a(N1624), .O(N1819) );
inv1 gate368( .a(N1619), .O(N1820) );
inv1 gate369( .a(N1615), .O(N1821) );
and4 gate370( .a(N496), .b(N224), .c(N36), .d(N1591), .O(N1822) );
and4 gate371( .a(N496), .b(N224), .c(N1591), .d(N486), .O(N1823) );
buf1 gate372( .a(N1596), .O(N1824) );
inv1 gate373( .a(N1606), .O(N1827) );
and2 gate374( .a(N1600), .b(N537), .O(N1830) );
and2 gate375( .a(N1606), .b(N537), .O(N1831) );
and2 gate376( .a(N1619), .b(N246), .O(N1832) );
inv1 gate377( .a(N1596), .O(N1833) );
inv1 gate378( .a(N1600), .O(N1836) );
inv1 gate379( .a(N1606), .O(N1841) );
buf1 gate380( .a(N1612), .O(N1848) );
buf1 gate381( .a(N1615), .O(N1852) );
buf1 gate382( .a(N1619), .O(N1856) );
buf1 gate383( .a(N1624), .O(N1863) );
buf1 gate384( .a(N1628), .O(N1870) );
buf1 gate385( .a(N1631), .O(N1875) );
buf1 gate386( .a(N1634), .O(N1880) );
nand2 gate387( .a(N727), .b(N1651), .O(N1885) );
nand2 gate388( .a(N730), .b(N1656), .O(N1888) );
buf1 gate389( .a(N1686), .O(N1891) );
and2 gate390( .a(N1637), .b(N425), .O(N1894) );
inv1 gate391( .a(N1642), .O(N1897) );
and3 gate392( .a(N1496), .b(N1133), .c(N1776), .O(N1908) );
and3 gate393( .a(N1129), .b(N1499), .c(N1777), .O(N1909) );
and2 gate394( .a(N1600), .b(N637), .O(N1910) );
and2 gate395( .a(N1606), .b(N637), .O(N1911) );
and2 gate396( .a(N1612), .b(N637), .O(N1912) );
and2 gate397( .a(N1615), .b(N637), .O(N1913) );
and2 gate398( .a(N1619), .b(N643), .O(N1914) );
and2 gate399( .a(N1624), .b(N643), .O(N1915) );
and2 gate400( .a(N1628), .b(N643), .O(N1916) );
and2 gate401( .a(N1631), .b(N643), .O(N1917) );
and2 gate402( .a(N1634), .b(N643), .O(N1918) );
inv1 gate403( .a(N1708), .O(N1919) );
and2 gate404( .a(N1676), .b(N693), .O(N1928) );
and2 gate405( .a(N1681), .b(N693), .O(N1929) );
and2 gate406( .a(N1686), .b(N693), .O(N1930) );
and2 gate407( .a(N1690), .b(N693), .O(N1931) );
and2 gate408( .a(N1637), .b(N699), .O(N1932) );
and2 gate409( .a(N1642), .b(N699), .O(N1933) );
and2 gate410( .a(N1647), .b(N699), .O(N1934) );
and2 gate411( .a(N1651), .b(N699), .O(N1935) );
buf1 gate412( .a(N1600), .O(N1936) );
nand2 gate413( .a(N1216), .b(N1808), .O(N1939) );
nand2 gate414( .a(N1585), .b(N1810), .O(N1940) );

  xor2  gate1564(.a(N1811), .b(N1582), .O(gate415inter0));
  nand2 gate1565(.a(gate415inter0), .b(s_42), .O(gate415inter1));
  and2  gate1566(.a(N1811), .b(N1582), .O(gate415inter2));
  inv1  gate1567(.a(s_42), .O(gate415inter3));
  inv1  gate1568(.a(s_43), .O(gate415inter4));
  nand2 gate1569(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1570(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1571(.a(N1582), .O(gate415inter7));
  inv1  gate1572(.a(N1811), .O(gate415inter8));
  nand2 gate1573(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1574(.a(s_43), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1575(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1576(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1577(.a(gate415inter12), .b(gate415inter1), .O(N1941));
buf1 gate416( .a(N1676), .O(N1942) );
buf1 gate417( .a(N1686), .O(N1945) );
buf1 gate418( .a(N1681), .O(N1948) );
buf1 gate419( .a(N1637), .O(N1951) );
buf1 gate420( .a(N1690), .O(N1954) );
buf1 gate421( .a(N1647), .O(N1957) );
buf1 gate422( .a(N1642), .O(N1960) );
buf1 gate423( .a(N1656), .O(N1963) );
buf1 gate424( .a(N1651), .O(N1966) );
or2 gate425( .a(N533), .b(N1815), .O(N1969) );
inv1 gate426( .a(N1822), .O(N1970) );
inv1 gate427( .a(N1823), .O(N1971) );
buf1 gate428( .a(N1848), .O(N2010) );
buf1 gate429( .a(N1852), .O(N2012) );
buf1 gate430( .a(N1856), .O(N2014) );
buf1 gate431( .a(N1863), .O(N2016) );
buf1 gate432( .a(N1870), .O(N2018) );
buf1 gate433( .a(N1875), .O(N2020) );
buf1 gate434( .a(N1880), .O(N2022) );
inv1 gate435( .a(N1778), .O(N2028) );
inv1 gate436( .a(N1781), .O(N2029) );
nor2 gate437( .a(N1908), .b(N1784), .O(N2030) );
nor2 gate438( .a(N1909), .b(N1785), .O(N2031) );
and3 gate439( .a(N1506), .b(N1502), .c(N1778), .O(N2032) );
and3 gate440( .a(N1773), .b(N1770), .c(N1781), .O(N2033) );
or2 gate441( .a(N1571), .b(N1935), .O(N2034) );
inv1 gate442( .a(N1801), .O(N2040) );
inv1 gate443( .a(N1804), .O(N2041) );
and3 gate444( .a(N1557), .b(N1553), .c(N1801), .O(N2042) );
and3 gate445( .a(N1798), .b(N1795), .c(N1804), .O(N2043) );
nand2 gate446( .a(N1939), .b(N1809), .O(N2046) );
nand2 gate447( .a(N1940), .b(N1941), .O(N2049) );
or2 gate448( .a(N1544), .b(N1910), .O(N2052) );
or2 gate449( .a(N1545), .b(N1911), .O(N2055) );
or2 gate450( .a(N1546), .b(N1912), .O(N2058) );
or2 gate451( .a(N1547), .b(N1913), .O(N2061) );
or2 gate452( .a(N1548), .b(N1914), .O(N2064) );
or2 gate453( .a(N1549), .b(N1915), .O(N2067) );
or2 gate454( .a(N1550), .b(N1916), .O(N2070) );
or2 gate455( .a(N1551), .b(N1917), .O(N2073) );
or2 gate456( .a(N1552), .b(N1918), .O(N2076) );
or2 gate457( .a(N1564), .b(N1928), .O(N2079) );
or2 gate458( .a(N1565), .b(N1929), .O(N2095) );
or2 gate459( .a(N1566), .b(N1930), .O(N2098) );
or2 gate460( .a(N1567), .b(N1931), .O(N2101) );
or2 gate461( .a(N1568), .b(N1932), .O(N2104) );
or2 gate462( .a(N1569), .b(N1933), .O(N2107) );
or2 gate463( .a(N1570), .b(N1934), .O(N2110) );
and3 gate464( .a(N1897), .b(N1894), .c(N40), .O(N2113) );
inv1 gate465( .a(N1894), .O(N2119) );
nand2 gate466( .a(N408), .b(N1827), .O(N2120) );
and2 gate467( .a(N1824), .b(N537), .O(N2125) );
and2 gate468( .a(N1852), .b(N246), .O(N2126) );
and2 gate469( .a(N1848), .b(N537), .O(N2127) );
inv1 gate470( .a(N1848), .O(N2128) );
inv1 gate471( .a(N1852), .O(N2135) );
inv1 gate472( .a(N1863), .O(N2141) );
inv1 gate473( .a(N1870), .O(N2144) );
inv1 gate474( .a(N1875), .O(N2147) );
inv1 gate475( .a(N1880), .O(N2150) );
and2 gate476( .a(N727), .b(N1885), .O(N2153) );
and2 gate477( .a(N1885), .b(N1651), .O(N2154) );
and2 gate478( .a(N730), .b(N1888), .O(N2155) );
and2 gate479( .a(N1888), .b(N1656), .O(N2156) );
and3 gate480( .a(N1770), .b(N1506), .c(N2028), .O(N2157) );
and3 gate481( .a(N1502), .b(N1773), .c(N2029), .O(N2158) );
inv1 gate482( .a(N1942), .O(N2171) );

  xor2  gate1718(.a(N1919), .b(N1942), .O(gate483inter0));
  nand2 gate1719(.a(gate483inter0), .b(s_64), .O(gate483inter1));
  and2  gate1720(.a(N1919), .b(N1942), .O(gate483inter2));
  inv1  gate1721(.a(s_64), .O(gate483inter3));
  inv1  gate1722(.a(s_65), .O(gate483inter4));
  nand2 gate1723(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1724(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1725(.a(N1942), .O(gate483inter7));
  inv1  gate1726(.a(N1919), .O(gate483inter8));
  nand2 gate1727(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1728(.a(s_65), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1729(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1730(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1731(.a(gate483inter12), .b(gate483inter1), .O(N2172));
inv1 gate484( .a(N1945), .O(N2173) );
inv1 gate485( .a(N1948), .O(N2174) );
inv1 gate486( .a(N1951), .O(N2175) );
inv1 gate487( .a(N1954), .O(N2176) );
and3 gate488( .a(N1795), .b(N1557), .c(N2040), .O(N2177) );
and3 gate489( .a(N1553), .b(N1798), .c(N2041), .O(N2178) );
buf1 gate490( .a(N1836), .O(N2185) );
buf1 gate491( .a(N1833), .O(N2188) );
buf1 gate492( .a(N1841), .O(N2191) );
inv1 gate493( .a(N1856), .O(N2194) );
inv1 gate494( .a(N1827), .O(N2197) );
inv1 gate495( .a(N1936), .O(N2200) );
buf1 gate496( .a(N1836), .O(N2201) );
buf1 gate497( .a(N1833), .O(N2204) );
buf1 gate498( .a(N1841), .O(N2207) );
buf1 gate499( .a(N1824), .O(N2210) );
buf1 gate500( .a(N1841), .O(N2213) );
buf1 gate501( .a(N1841), .O(N2216) );
nand2 gate502( .a(N2031), .b(N2030), .O(N2219) );
inv1 gate503( .a(N1957), .O(N2234) );
inv1 gate504( .a(N1960), .O(N2235) );
inv1 gate505( .a(N1963), .O(N2236) );
inv1 gate506( .a(N1966), .O(N2237) );
and3 gate507( .a(N40), .b(N1897), .c(N2119), .O(N2250) );
or2 gate508( .a(N1831), .b(N2126), .O(N2266) );
or2 gate509( .a(N2127), .b(N1832), .O(N2269) );
or2 gate510( .a(N2153), .b(N2154), .O(N2291) );
or2 gate511( .a(N2155), .b(N2156), .O(N2294) );
nor2 gate512( .a(N2157), .b(N2032), .O(N2297) );
nor2 gate513( .a(N2158), .b(N2033), .O(N2298) );
inv1 gate514( .a(N2046), .O(N2300) );
inv1 gate515( .a(N2049), .O(N2301) );
nand2 gate516( .a(N2052), .b(N1519), .O(N2302) );
inv1 gate517( .a(N2052), .O(N2303) );
nand2 gate518( .a(N2055), .b(N1520), .O(N2304) );
inv1 gate519( .a(N2055), .O(N2305) );
nand2 gate520( .a(N2058), .b(N1521), .O(N2306) );
inv1 gate521( .a(N2058), .O(N2307) );
nand2 gate522( .a(N2061), .b(N1522), .O(N2308) );
inv1 gate523( .a(N2061), .O(N2309) );
nand2 gate524( .a(N2064), .b(N1523), .O(N2310) );
inv1 gate525( .a(N2064), .O(N2311) );
nand2 gate526( .a(N2067), .b(N1524), .O(N2312) );
inv1 gate527( .a(N2067), .O(N2313) );
nand2 gate528( .a(N2070), .b(N1525), .O(N2314) );
inv1 gate529( .a(N2070), .O(N2315) );
nand2 gate530( .a(N2073), .b(N1526), .O(N2316) );
inv1 gate531( .a(N2073), .O(N2317) );

  xor2  gate1466(.a(N1527), .b(N2076), .O(gate532inter0));
  nand2 gate1467(.a(gate532inter0), .b(s_28), .O(gate532inter1));
  and2  gate1468(.a(N1527), .b(N2076), .O(gate532inter2));
  inv1  gate1469(.a(s_28), .O(gate532inter3));
  inv1  gate1470(.a(s_29), .O(gate532inter4));
  nand2 gate1471(.a(gate532inter4), .b(gate532inter3), .O(gate532inter5));
  nor2  gate1472(.a(gate532inter5), .b(gate532inter2), .O(gate532inter6));
  inv1  gate1473(.a(N2076), .O(gate532inter7));
  inv1  gate1474(.a(N1527), .O(gate532inter8));
  nand2 gate1475(.a(gate532inter8), .b(gate532inter7), .O(gate532inter9));
  nand2 gate1476(.a(s_29), .b(gate532inter3), .O(gate532inter10));
  nor2  gate1477(.a(gate532inter10), .b(gate532inter9), .O(gate532inter11));
  nor2  gate1478(.a(gate532inter11), .b(gate532inter6), .O(gate532inter12));
  nand2 gate1479(.a(gate532inter12), .b(gate532inter1), .O(N2318));
inv1 gate533( .a(N2076), .O(N2319) );

  xor2  gate1928(.a(N1528), .b(N2079), .O(gate534inter0));
  nand2 gate1929(.a(gate534inter0), .b(s_94), .O(gate534inter1));
  and2  gate1930(.a(N1528), .b(N2079), .O(gate534inter2));
  inv1  gate1931(.a(s_94), .O(gate534inter3));
  inv1  gate1932(.a(s_95), .O(gate534inter4));
  nand2 gate1933(.a(gate534inter4), .b(gate534inter3), .O(gate534inter5));
  nor2  gate1934(.a(gate534inter5), .b(gate534inter2), .O(gate534inter6));
  inv1  gate1935(.a(N2079), .O(gate534inter7));
  inv1  gate1936(.a(N1528), .O(gate534inter8));
  nand2 gate1937(.a(gate534inter8), .b(gate534inter7), .O(gate534inter9));
  nand2 gate1938(.a(s_95), .b(gate534inter3), .O(gate534inter10));
  nor2  gate1939(.a(gate534inter10), .b(gate534inter9), .O(gate534inter11));
  nor2  gate1940(.a(gate534inter11), .b(gate534inter6), .O(gate534inter12));
  nand2 gate1941(.a(gate534inter12), .b(gate534inter1), .O(N2320));
inv1 gate535( .a(N2079), .O(N2321) );

  xor2  gate1914(.a(N2171), .b(N1708), .O(gate536inter0));
  nand2 gate1915(.a(gate536inter0), .b(s_92), .O(gate536inter1));
  and2  gate1916(.a(N2171), .b(N1708), .O(gate536inter2));
  inv1  gate1917(.a(s_92), .O(gate536inter3));
  inv1  gate1918(.a(s_93), .O(gate536inter4));
  nand2 gate1919(.a(gate536inter4), .b(gate536inter3), .O(gate536inter5));
  nor2  gate1920(.a(gate536inter5), .b(gate536inter2), .O(gate536inter6));
  inv1  gate1921(.a(N1708), .O(gate536inter7));
  inv1  gate1922(.a(N2171), .O(gate536inter8));
  nand2 gate1923(.a(gate536inter8), .b(gate536inter7), .O(gate536inter9));
  nand2 gate1924(.a(s_93), .b(gate536inter3), .O(gate536inter10));
  nor2  gate1925(.a(gate536inter10), .b(gate536inter9), .O(gate536inter11));
  nor2  gate1926(.a(gate536inter11), .b(gate536inter6), .O(gate536inter12));
  nand2 gate1927(.a(gate536inter12), .b(gate536inter1), .O(N2322));
nand2 gate537( .a(N1948), .b(N2173), .O(N2323) );

  xor2  gate1648(.a(N2174), .b(N1945), .O(gate538inter0));
  nand2 gate1649(.a(gate538inter0), .b(s_54), .O(gate538inter1));
  and2  gate1650(.a(N2174), .b(N1945), .O(gate538inter2));
  inv1  gate1651(.a(s_54), .O(gate538inter3));
  inv1  gate1652(.a(s_55), .O(gate538inter4));
  nand2 gate1653(.a(gate538inter4), .b(gate538inter3), .O(gate538inter5));
  nor2  gate1654(.a(gate538inter5), .b(gate538inter2), .O(gate538inter6));
  inv1  gate1655(.a(N1945), .O(gate538inter7));
  inv1  gate1656(.a(N2174), .O(gate538inter8));
  nand2 gate1657(.a(gate538inter8), .b(gate538inter7), .O(gate538inter9));
  nand2 gate1658(.a(s_55), .b(gate538inter3), .O(gate538inter10));
  nor2  gate1659(.a(gate538inter10), .b(gate538inter9), .O(gate538inter11));
  nor2  gate1660(.a(gate538inter11), .b(gate538inter6), .O(gate538inter12));
  nand2 gate1661(.a(gate538inter12), .b(gate538inter1), .O(N2324));
nand2 gate539( .a(N1954), .b(N2175), .O(N2325) );
nand2 gate540( .a(N1951), .b(N2176), .O(N2326) );
nor2 gate541( .a(N2177), .b(N2042), .O(N2327) );
nor2 gate542( .a(N2178), .b(N2043), .O(N2328) );
nand2 gate543( .a(N2095), .b(N1572), .O(N2329) );
inv1 gate544( .a(N2095), .O(N2330) );
nand2 gate545( .a(N2098), .b(N1573), .O(N2331) );
inv1 gate546( .a(N2098), .O(N2332) );
nand2 gate547( .a(N2101), .b(N1574), .O(N2333) );
inv1 gate548( .a(N2101), .O(N2334) );
nand2 gate549( .a(N2104), .b(N1575), .O(N2335) );
inv1 gate550( .a(N2104), .O(N2336) );
nand2 gate551( .a(N2107), .b(N1576), .O(N2337) );
inv1 gate552( .a(N2107), .O(N2338) );
nand2 gate553( .a(N2110), .b(N1577), .O(N2339) );
inv1 gate554( .a(N2110), .O(N2340) );

  xor2  gate1550(.a(N2234), .b(N1960), .O(gate555inter0));
  nand2 gate1551(.a(gate555inter0), .b(s_40), .O(gate555inter1));
  and2  gate1552(.a(N2234), .b(N1960), .O(gate555inter2));
  inv1  gate1553(.a(s_40), .O(gate555inter3));
  inv1  gate1554(.a(s_41), .O(gate555inter4));
  nand2 gate1555(.a(gate555inter4), .b(gate555inter3), .O(gate555inter5));
  nor2  gate1556(.a(gate555inter5), .b(gate555inter2), .O(gate555inter6));
  inv1  gate1557(.a(N1960), .O(gate555inter7));
  inv1  gate1558(.a(N2234), .O(gate555inter8));
  nand2 gate1559(.a(gate555inter8), .b(gate555inter7), .O(gate555inter9));
  nand2 gate1560(.a(s_41), .b(gate555inter3), .O(gate555inter10));
  nor2  gate1561(.a(gate555inter10), .b(gate555inter9), .O(gate555inter11));
  nor2  gate1562(.a(gate555inter11), .b(gate555inter6), .O(gate555inter12));
  nand2 gate1563(.a(gate555inter12), .b(gate555inter1), .O(N2354));
nand2 gate556( .a(N1957), .b(N2235), .O(N2355) );
nand2 gate557( .a(N1966), .b(N2236), .O(N2356) );

  xor2  gate1998(.a(N2237), .b(N1963), .O(gate558inter0));
  nand2 gate1999(.a(gate558inter0), .b(s_104), .O(gate558inter1));
  and2  gate2000(.a(N2237), .b(N1963), .O(gate558inter2));
  inv1  gate2001(.a(s_104), .O(gate558inter3));
  inv1  gate2002(.a(s_105), .O(gate558inter4));
  nand2 gate2003(.a(gate558inter4), .b(gate558inter3), .O(gate558inter5));
  nor2  gate2004(.a(gate558inter5), .b(gate558inter2), .O(gate558inter6));
  inv1  gate2005(.a(N1963), .O(gate558inter7));
  inv1  gate2006(.a(N2237), .O(gate558inter8));
  nand2 gate2007(.a(gate558inter8), .b(gate558inter7), .O(gate558inter9));
  nand2 gate2008(.a(s_105), .b(gate558inter3), .O(gate558inter10));
  nor2  gate2009(.a(gate558inter10), .b(gate558inter9), .O(gate558inter11));
  nor2  gate2010(.a(gate558inter11), .b(gate558inter6), .O(gate558inter12));
  nand2 gate2011(.a(gate558inter12), .b(gate558inter1), .O(N2357));
and2 gate559( .a(N2120), .b(N533), .O(N2358) );
inv1 gate560( .a(N2113), .O(N2359) );
inv1 gate561( .a(N2185), .O(N2364) );
inv1 gate562( .a(N2188), .O(N2365) );
inv1 gate563( .a(N2191), .O(N2366) );
inv1 gate564( .a(N2194), .O(N2367) );
buf1 gate565( .a(N2120), .O(N2368) );
inv1 gate566( .a(N2201), .O(N2372) );
inv1 gate567( .a(N2204), .O(N2373) );
inv1 gate568( .a(N2207), .O(N2374) );
inv1 gate569( .a(N2210), .O(N2375) );
inv1 gate570( .a(N2213), .O(N2376) );
inv1 gate571( .a(N2113), .O(N2377) );
buf1 gate572( .a(N2113), .O(N2382) );
and2 gate573( .a(N2120), .b(N246), .O(N2386) );
buf1 gate574( .a(N2266), .O(N2387) );
buf1 gate575( .a(N2266), .O(N2388) );
buf1 gate576( .a(N2269), .O(N2389) );
buf1 gate577( .a(N2269), .O(N2390) );
buf1 gate578( .a(N2113), .O(N2391) );
inv1 gate579( .a(N2113), .O(N2395) );
nand2 gate580( .a(N2219), .b(N2300), .O(N2400) );
inv1 gate581( .a(N2216), .O(N2403) );
inv1 gate582( .a(N2219), .O(N2406) );

  xor2  gate1592(.a(N2303), .b(N1219), .O(gate583inter0));
  nand2 gate1593(.a(gate583inter0), .b(s_46), .O(gate583inter1));
  and2  gate1594(.a(N2303), .b(N1219), .O(gate583inter2));
  inv1  gate1595(.a(s_46), .O(gate583inter3));
  inv1  gate1596(.a(s_47), .O(gate583inter4));
  nand2 gate1597(.a(gate583inter4), .b(gate583inter3), .O(gate583inter5));
  nor2  gate1598(.a(gate583inter5), .b(gate583inter2), .O(gate583inter6));
  inv1  gate1599(.a(N1219), .O(gate583inter7));
  inv1  gate1600(.a(N2303), .O(gate583inter8));
  nand2 gate1601(.a(gate583inter8), .b(gate583inter7), .O(gate583inter9));
  nand2 gate1602(.a(s_47), .b(gate583inter3), .O(gate583inter10));
  nor2  gate1603(.a(gate583inter10), .b(gate583inter9), .O(gate583inter11));
  nor2  gate1604(.a(gate583inter11), .b(gate583inter6), .O(gate583inter12));
  nand2 gate1605(.a(gate583inter12), .b(gate583inter1), .O(N2407));
nand2 gate584( .a(N1222), .b(N2305), .O(N2408) );
nand2 gate585( .a(N1225), .b(N2307), .O(N2409) );

  xor2  gate2012(.a(N2309), .b(N1228), .O(gate586inter0));
  nand2 gate2013(.a(gate586inter0), .b(s_106), .O(gate586inter1));
  and2  gate2014(.a(N2309), .b(N1228), .O(gate586inter2));
  inv1  gate2015(.a(s_106), .O(gate586inter3));
  inv1  gate2016(.a(s_107), .O(gate586inter4));
  nand2 gate2017(.a(gate586inter4), .b(gate586inter3), .O(gate586inter5));
  nor2  gate2018(.a(gate586inter5), .b(gate586inter2), .O(gate586inter6));
  inv1  gate2019(.a(N1228), .O(gate586inter7));
  inv1  gate2020(.a(N2309), .O(gate586inter8));
  nand2 gate2021(.a(gate586inter8), .b(gate586inter7), .O(gate586inter9));
  nand2 gate2022(.a(s_107), .b(gate586inter3), .O(gate586inter10));
  nor2  gate2023(.a(gate586inter10), .b(gate586inter9), .O(gate586inter11));
  nor2  gate2024(.a(gate586inter11), .b(gate586inter6), .O(gate586inter12));
  nand2 gate2025(.a(gate586inter12), .b(gate586inter1), .O(N2410));

  xor2  gate1424(.a(N2311), .b(N1231), .O(gate587inter0));
  nand2 gate1425(.a(gate587inter0), .b(s_22), .O(gate587inter1));
  and2  gate1426(.a(N2311), .b(N1231), .O(gate587inter2));
  inv1  gate1427(.a(s_22), .O(gate587inter3));
  inv1  gate1428(.a(s_23), .O(gate587inter4));
  nand2 gate1429(.a(gate587inter4), .b(gate587inter3), .O(gate587inter5));
  nor2  gate1430(.a(gate587inter5), .b(gate587inter2), .O(gate587inter6));
  inv1  gate1431(.a(N1231), .O(gate587inter7));
  inv1  gate1432(.a(N2311), .O(gate587inter8));
  nand2 gate1433(.a(gate587inter8), .b(gate587inter7), .O(gate587inter9));
  nand2 gate1434(.a(s_23), .b(gate587inter3), .O(gate587inter10));
  nor2  gate1435(.a(gate587inter10), .b(gate587inter9), .O(gate587inter11));
  nor2  gate1436(.a(gate587inter11), .b(gate587inter6), .O(gate587inter12));
  nand2 gate1437(.a(gate587inter12), .b(gate587inter1), .O(N2411));
nand2 gate588( .a(N1234), .b(N2313), .O(N2412) );
nand2 gate589( .a(N1237), .b(N2315), .O(N2413) );
nand2 gate590( .a(N1240), .b(N2317), .O(N2414) );

  xor2  gate1298(.a(N2319), .b(N1243), .O(gate591inter0));
  nand2 gate1299(.a(gate591inter0), .b(s_4), .O(gate591inter1));
  and2  gate1300(.a(N2319), .b(N1243), .O(gate591inter2));
  inv1  gate1301(.a(s_4), .O(gate591inter3));
  inv1  gate1302(.a(s_5), .O(gate591inter4));
  nand2 gate1303(.a(gate591inter4), .b(gate591inter3), .O(gate591inter5));
  nor2  gate1304(.a(gate591inter5), .b(gate591inter2), .O(gate591inter6));
  inv1  gate1305(.a(N1243), .O(gate591inter7));
  inv1  gate1306(.a(N2319), .O(gate591inter8));
  nand2 gate1307(.a(gate591inter8), .b(gate591inter7), .O(gate591inter9));
  nand2 gate1308(.a(s_5), .b(gate591inter3), .O(gate591inter10));
  nor2  gate1309(.a(gate591inter10), .b(gate591inter9), .O(gate591inter11));
  nor2  gate1310(.a(gate591inter11), .b(gate591inter6), .O(gate591inter12));
  nand2 gate1311(.a(gate591inter12), .b(gate591inter1), .O(N2415));
nand2 gate592( .a(N1246), .b(N2321), .O(N2416) );
nand2 gate593( .a(N2322), .b(N2172), .O(N2417) );
nand2 gate594( .a(N2323), .b(N2324), .O(N2421) );
nand2 gate595( .a(N2325), .b(N2326), .O(N2425) );
nand2 gate596( .a(N1251), .b(N2330), .O(N2428) );
nand2 gate597( .a(N1254), .b(N2332), .O(N2429) );
nand2 gate598( .a(N1257), .b(N2334), .O(N2430) );
nand2 gate599( .a(N1260), .b(N2336), .O(N2431) );
nand2 gate600( .a(N1263), .b(N2338), .O(N2432) );
nand2 gate601( .a(N1266), .b(N2340), .O(N2433) );
buf1 gate602( .a(N2128), .O(N2434) );
buf1 gate603( .a(N2135), .O(N2437) );
buf1 gate604( .a(N2144), .O(N2440) );
buf1 gate605( .a(N2141), .O(N2443) );
buf1 gate606( .a(N2150), .O(N2446) );
buf1 gate607( .a(N2147), .O(N2449) );
inv1 gate608( .a(N2197), .O(N2452) );

  xor2  gate1956(.a(N2200), .b(N2197), .O(gate609inter0));
  nand2 gate1957(.a(gate609inter0), .b(s_98), .O(gate609inter1));
  and2  gate1958(.a(N2200), .b(N2197), .O(gate609inter2));
  inv1  gate1959(.a(s_98), .O(gate609inter3));
  inv1  gate1960(.a(s_99), .O(gate609inter4));
  nand2 gate1961(.a(gate609inter4), .b(gate609inter3), .O(gate609inter5));
  nor2  gate1962(.a(gate609inter5), .b(gate609inter2), .O(gate609inter6));
  inv1  gate1963(.a(N2197), .O(gate609inter7));
  inv1  gate1964(.a(N2200), .O(gate609inter8));
  nand2 gate1965(.a(gate609inter8), .b(gate609inter7), .O(gate609inter9));
  nand2 gate1966(.a(s_99), .b(gate609inter3), .O(gate609inter10));
  nor2  gate1967(.a(gate609inter10), .b(gate609inter9), .O(gate609inter11));
  nor2  gate1968(.a(gate609inter11), .b(gate609inter6), .O(gate609inter12));
  nand2 gate1969(.a(gate609inter12), .b(gate609inter1), .O(N2453));
buf1 gate610( .a(N2128), .O(N2454) );
buf1 gate611( .a(N2144), .O(N2457) );
buf1 gate612( .a(N2141), .O(N2460) );
buf1 gate613( .a(N2150), .O(N2463) );
buf1 gate614( .a(N2147), .O(N2466) );
inv1 gate615( .a(N2120), .O(N2469) );
buf1 gate616( .a(N2128), .O(N2472) );
buf1 gate617( .a(N2135), .O(N2475) );
buf1 gate618( .a(N2128), .O(N2478) );
buf1 gate619( .a(N2135), .O(N2481) );
nand2 gate620( .a(N2298), .b(N2297), .O(N2484) );
nand2 gate621( .a(N2356), .b(N2357), .O(N2487) );
nand2 gate622( .a(N2354), .b(N2355), .O(N2490) );
nand2 gate623( .a(N2328), .b(N2327), .O(N2493) );
or2 gate624( .a(N2358), .b(N1814), .O(N2496) );
nand2 gate625( .a(N2188), .b(N2364), .O(N2503) );
nand2 gate626( .a(N2185), .b(N2365), .O(N2504) );
nand2 gate627( .a(N2204), .b(N2372), .O(N2510) );
nand2 gate628( .a(N2201), .b(N2373), .O(N2511) );
or2 gate629( .a(N1830), .b(N2386), .O(N2521) );
nand2 gate630( .a(N2046), .b(N2406), .O(N2528) );
inv1 gate631( .a(N2291), .O(N2531) );
inv1 gate632( .a(N2294), .O(N2534) );
buf1 gate633( .a(N2250), .O(N2537) );
buf1 gate634( .a(N2250), .O(N2540) );
nand2 gate635( .a(N2302), .b(N2407), .O(N2544) );
nand2 gate636( .a(N2304), .b(N2408), .O(N2545) );
nand2 gate637( .a(N2306), .b(N2409), .O(N2546) );

  xor2  gate1844(.a(N2410), .b(N2308), .O(gate638inter0));
  nand2 gate1845(.a(gate638inter0), .b(s_82), .O(gate638inter1));
  and2  gate1846(.a(N2410), .b(N2308), .O(gate638inter2));
  inv1  gate1847(.a(s_82), .O(gate638inter3));
  inv1  gate1848(.a(s_83), .O(gate638inter4));
  nand2 gate1849(.a(gate638inter4), .b(gate638inter3), .O(gate638inter5));
  nor2  gate1850(.a(gate638inter5), .b(gate638inter2), .O(gate638inter6));
  inv1  gate1851(.a(N2308), .O(gate638inter7));
  inv1  gate1852(.a(N2410), .O(gate638inter8));
  nand2 gate1853(.a(gate638inter8), .b(gate638inter7), .O(gate638inter9));
  nand2 gate1854(.a(s_83), .b(gate638inter3), .O(gate638inter10));
  nor2  gate1855(.a(gate638inter10), .b(gate638inter9), .O(gate638inter11));
  nor2  gate1856(.a(gate638inter11), .b(gate638inter6), .O(gate638inter12));
  nand2 gate1857(.a(gate638inter12), .b(gate638inter1), .O(N2547));
nand2 gate639( .a(N2310), .b(N2411), .O(N2548) );
nand2 gate640( .a(N2312), .b(N2412), .O(N2549) );

  xor2  gate1578(.a(N2413), .b(N2314), .O(gate641inter0));
  nand2 gate1579(.a(gate641inter0), .b(s_44), .O(gate641inter1));
  and2  gate1580(.a(N2413), .b(N2314), .O(gate641inter2));
  inv1  gate1581(.a(s_44), .O(gate641inter3));
  inv1  gate1582(.a(s_45), .O(gate641inter4));
  nand2 gate1583(.a(gate641inter4), .b(gate641inter3), .O(gate641inter5));
  nor2  gate1584(.a(gate641inter5), .b(gate641inter2), .O(gate641inter6));
  inv1  gate1585(.a(N2314), .O(gate641inter7));
  inv1  gate1586(.a(N2413), .O(gate641inter8));
  nand2 gate1587(.a(gate641inter8), .b(gate641inter7), .O(gate641inter9));
  nand2 gate1588(.a(s_45), .b(gate641inter3), .O(gate641inter10));
  nor2  gate1589(.a(gate641inter10), .b(gate641inter9), .O(gate641inter11));
  nor2  gate1590(.a(gate641inter11), .b(gate641inter6), .O(gate641inter12));
  nand2 gate1591(.a(gate641inter12), .b(gate641inter1), .O(N2550));
nand2 gate642( .a(N2316), .b(N2414), .O(N2551) );
nand2 gate643( .a(N2318), .b(N2415), .O(N2552) );

  xor2  gate1872(.a(N2416), .b(N2320), .O(gate644inter0));
  nand2 gate1873(.a(gate644inter0), .b(s_86), .O(gate644inter1));
  and2  gate1874(.a(N2416), .b(N2320), .O(gate644inter2));
  inv1  gate1875(.a(s_86), .O(gate644inter3));
  inv1  gate1876(.a(s_87), .O(gate644inter4));
  nand2 gate1877(.a(gate644inter4), .b(gate644inter3), .O(gate644inter5));
  nor2  gate1878(.a(gate644inter5), .b(gate644inter2), .O(gate644inter6));
  inv1  gate1879(.a(N2320), .O(gate644inter7));
  inv1  gate1880(.a(N2416), .O(gate644inter8));
  nand2 gate1881(.a(gate644inter8), .b(gate644inter7), .O(gate644inter9));
  nand2 gate1882(.a(s_87), .b(gate644inter3), .O(gate644inter10));
  nor2  gate1883(.a(gate644inter10), .b(gate644inter9), .O(gate644inter11));
  nor2  gate1884(.a(gate644inter11), .b(gate644inter6), .O(gate644inter12));
  nand2 gate1885(.a(gate644inter12), .b(gate644inter1), .O(N2553));
nand2 gate645( .a(N2329), .b(N2428), .O(N2563) );

  xor2  gate1662(.a(N2429), .b(N2331), .O(gate646inter0));
  nand2 gate1663(.a(gate646inter0), .b(s_56), .O(gate646inter1));
  and2  gate1664(.a(N2429), .b(N2331), .O(gate646inter2));
  inv1  gate1665(.a(s_56), .O(gate646inter3));
  inv1  gate1666(.a(s_57), .O(gate646inter4));
  nand2 gate1667(.a(gate646inter4), .b(gate646inter3), .O(gate646inter5));
  nor2  gate1668(.a(gate646inter5), .b(gate646inter2), .O(gate646inter6));
  inv1  gate1669(.a(N2331), .O(gate646inter7));
  inv1  gate1670(.a(N2429), .O(gate646inter8));
  nand2 gate1671(.a(gate646inter8), .b(gate646inter7), .O(gate646inter9));
  nand2 gate1672(.a(s_57), .b(gate646inter3), .O(gate646inter10));
  nor2  gate1673(.a(gate646inter10), .b(gate646inter9), .O(gate646inter11));
  nor2  gate1674(.a(gate646inter11), .b(gate646inter6), .O(gate646inter12));
  nand2 gate1675(.a(gate646inter12), .b(gate646inter1), .O(N2564));

  xor2  gate1732(.a(N2430), .b(N2333), .O(gate647inter0));
  nand2 gate1733(.a(gate647inter0), .b(s_66), .O(gate647inter1));
  and2  gate1734(.a(N2430), .b(N2333), .O(gate647inter2));
  inv1  gate1735(.a(s_66), .O(gate647inter3));
  inv1  gate1736(.a(s_67), .O(gate647inter4));
  nand2 gate1737(.a(gate647inter4), .b(gate647inter3), .O(gate647inter5));
  nor2  gate1738(.a(gate647inter5), .b(gate647inter2), .O(gate647inter6));
  inv1  gate1739(.a(N2333), .O(gate647inter7));
  inv1  gate1740(.a(N2430), .O(gate647inter8));
  nand2 gate1741(.a(gate647inter8), .b(gate647inter7), .O(gate647inter9));
  nand2 gate1742(.a(s_67), .b(gate647inter3), .O(gate647inter10));
  nor2  gate1743(.a(gate647inter10), .b(gate647inter9), .O(gate647inter11));
  nor2  gate1744(.a(gate647inter11), .b(gate647inter6), .O(gate647inter12));
  nand2 gate1745(.a(gate647inter12), .b(gate647inter1), .O(N2565));
nand2 gate648( .a(N2335), .b(N2431), .O(N2566) );
nand2 gate649( .a(N2337), .b(N2432), .O(N2567) );

  xor2  gate1396(.a(N2433), .b(N2339), .O(gate650inter0));
  nand2 gate1397(.a(gate650inter0), .b(s_18), .O(gate650inter1));
  and2  gate1398(.a(N2433), .b(N2339), .O(gate650inter2));
  inv1  gate1399(.a(s_18), .O(gate650inter3));
  inv1  gate1400(.a(s_19), .O(gate650inter4));
  nand2 gate1401(.a(gate650inter4), .b(gate650inter3), .O(gate650inter5));
  nor2  gate1402(.a(gate650inter5), .b(gate650inter2), .O(gate650inter6));
  inv1  gate1403(.a(N2339), .O(gate650inter7));
  inv1  gate1404(.a(N2433), .O(gate650inter8));
  nand2 gate1405(.a(gate650inter8), .b(gate650inter7), .O(gate650inter9));
  nand2 gate1406(.a(s_19), .b(gate650inter3), .O(gate650inter10));
  nor2  gate1407(.a(gate650inter10), .b(gate650inter9), .O(gate650inter11));
  nor2  gate1408(.a(gate650inter11), .b(gate650inter6), .O(gate650inter12));
  nand2 gate1409(.a(gate650inter12), .b(gate650inter1), .O(N2568));

  xor2  gate1382(.a(N2452), .b(N1936), .O(gate651inter0));
  nand2 gate1383(.a(gate651inter0), .b(s_16), .O(gate651inter1));
  and2  gate1384(.a(N2452), .b(N1936), .O(gate651inter2));
  inv1  gate1385(.a(s_16), .O(gate651inter3));
  inv1  gate1386(.a(s_17), .O(gate651inter4));
  nand2 gate1387(.a(gate651inter4), .b(gate651inter3), .O(gate651inter5));
  nor2  gate1388(.a(gate651inter5), .b(gate651inter2), .O(gate651inter6));
  inv1  gate1389(.a(N1936), .O(gate651inter7));
  inv1  gate1390(.a(N2452), .O(gate651inter8));
  nand2 gate1391(.a(gate651inter8), .b(gate651inter7), .O(gate651inter9));
  nand2 gate1392(.a(s_17), .b(gate651inter3), .O(gate651inter10));
  nor2  gate1393(.a(gate651inter10), .b(gate651inter9), .O(gate651inter11));
  nor2  gate1394(.a(gate651inter11), .b(gate651inter6), .O(gate651inter12));
  nand2 gate1395(.a(gate651inter12), .b(gate651inter1), .O(N2579));
buf1 gate652( .a(N2359), .O(N2603) );
and2 gate653( .a(N1880), .b(N2377), .O(N2607) );
and2 gate654( .a(N1676), .b(N2377), .O(N2608) );
and2 gate655( .a(N1681), .b(N2377), .O(N2609) );
and2 gate656( .a(N1891), .b(N2377), .O(N2610) );
and2 gate657( .a(N1856), .b(N2382), .O(N2611) );
and2 gate658( .a(N1863), .b(N2382), .O(N2612) );
nand2 gate659( .a(N2503), .b(N2504), .O(N2613) );
inv1 gate660( .a(N2434), .O(N2617) );
nand2 gate661( .a(N2434), .b(N2366), .O(N2618) );
nand2 gate662( .a(N2437), .b(N2367), .O(N2619) );
inv1 gate663( .a(N2437), .O(N2620) );
inv1 gate664( .a(N2368), .O(N2621) );
nand2 gate665( .a(N2510), .b(N2511), .O(N2624) );
inv1 gate666( .a(N2454), .O(N2628) );
nand2 gate667( .a(N2454), .b(N2374), .O(N2629) );
inv1 gate668( .a(N2472), .O(N2630) );
and2 gate669( .a(N1856), .b(N2391), .O(N2631) );
and2 gate670( .a(N1863), .b(N2391), .O(N2632) );
and2 gate671( .a(N1880), .b(N2395), .O(N2633) );
and2 gate672( .a(N1676), .b(N2395), .O(N2634) );
and2 gate673( .a(N1681), .b(N2395), .O(N2635) );
and2 gate674( .a(N1891), .b(N2395), .O(N2636) );
inv1 gate675( .a(N2382), .O(N2638) );
buf1 gate676( .a(N2521), .O(N2643) );
buf1 gate677( .a(N2521), .O(N2644) );
inv1 gate678( .a(N2475), .O(N2645) );
inv1 gate679( .a(N2391), .O(N2646) );
nand2 gate680( .a(N2528), .b(N2400), .O(N2652) );
inv1 gate681( .a(N2478), .O(N2655) );
inv1 gate682( .a(N2481), .O(N2656) );
buf1 gate683( .a(N2359), .O(N2659) );
inv1 gate684( .a(N2484), .O(N2663) );
nand2 gate685( .a(N2484), .b(N2301), .O(N2664) );
inv1 gate686( .a(N2553), .O(N2665) );
inv1 gate687( .a(N2552), .O(N2666) );
inv1 gate688( .a(N2551), .O(N2667) );
inv1 gate689( .a(N2550), .O(N2668) );
inv1 gate690( .a(N2549), .O(N2669) );
inv1 gate691( .a(N2548), .O(N2670) );
inv1 gate692( .a(N2547), .O(N2671) );
inv1 gate693( .a(N2546), .O(N2672) );
inv1 gate694( .a(N2545), .O(N2673) );
inv1 gate695( .a(N2544), .O(N2674) );
inv1 gate696( .a(N2568), .O(N2675) );
inv1 gate697( .a(N2567), .O(N2676) );
inv1 gate698( .a(N2566), .O(N2677) );
inv1 gate699( .a(N2565), .O(N2678) );
inv1 gate700( .a(N2564), .O(N2679) );
inv1 gate701( .a(N2563), .O(N2680) );
inv1 gate702( .a(N2417), .O(N2681) );
inv1 gate703( .a(N2421), .O(N2684) );
buf1 gate704( .a(N2425), .O(N2687) );
buf1 gate705( .a(N2425), .O(N2690) );
inv1 gate706( .a(N2493), .O(N2693) );
nand2 gate707( .a(N2493), .b(N1807), .O(N2694) );
inv1 gate708( .a(N2440), .O(N2695) );
inv1 gate709( .a(N2443), .O(N2696) );
inv1 gate710( .a(N2446), .O(N2697) );
inv1 gate711( .a(N2449), .O(N2698) );
inv1 gate712( .a(N2457), .O(N2699) );
inv1 gate713( .a(N2460), .O(N2700) );
inv1 gate714( .a(N2463), .O(N2701) );
inv1 gate715( .a(N2466), .O(N2702) );

  xor2  gate1354(.a(N2453), .b(N2579), .O(gate716inter0));
  nand2 gate1355(.a(gate716inter0), .b(s_12), .O(gate716inter1));
  and2  gate1356(.a(N2453), .b(N2579), .O(gate716inter2));
  inv1  gate1357(.a(s_12), .O(gate716inter3));
  inv1  gate1358(.a(s_13), .O(gate716inter4));
  nand2 gate1359(.a(gate716inter4), .b(gate716inter3), .O(gate716inter5));
  nor2  gate1360(.a(gate716inter5), .b(gate716inter2), .O(gate716inter6));
  inv1  gate1361(.a(N2579), .O(gate716inter7));
  inv1  gate1362(.a(N2453), .O(gate716inter8));
  nand2 gate1363(.a(gate716inter8), .b(gate716inter7), .O(gate716inter9));
  nand2 gate1364(.a(s_13), .b(gate716inter3), .O(gate716inter10));
  nor2  gate1365(.a(gate716inter10), .b(gate716inter9), .O(gate716inter11));
  nor2  gate1366(.a(gate716inter11), .b(gate716inter6), .O(gate716inter12));
  nand2 gate1367(.a(gate716inter12), .b(gate716inter1), .O(N2703));
inv1 gate717( .a(N2469), .O(N2706) );
inv1 gate718( .a(N2487), .O(N2707) );
inv1 gate719( .a(N2490), .O(N2708) );
and2 gate720( .a(N2294), .b(N2534), .O(N2709) );
and2 gate721( .a(N2291), .b(N2531), .O(N2710) );
nand2 gate722( .a(N2191), .b(N2617), .O(N2719) );
nand2 gate723( .a(N2194), .b(N2620), .O(N2720) );
nand2 gate724( .a(N2207), .b(N2628), .O(N2726) );
buf1 gate725( .a(N2537), .O(N2729) );
buf1 gate726( .a(N2537), .O(N2738) );
inv1 gate727( .a(N2652), .O(N2743) );
nand2 gate728( .a(N2049), .b(N2663), .O(N2747) );
and5 gate729( .a(N2665), .b(N2666), .c(N2667), .d(N2668), .e(N2669), .O(N2748) );
and5 gate730( .a(N2670), .b(N2671), .c(N2672), .d(N2673), .e(N2674), .O(N2749) );
and2 gate731( .a(N2034), .b(N2675), .O(N2750) );
and5 gate732( .a(N2676), .b(N2677), .c(N2678), .d(N2679), .e(N2680), .O(N2751) );
nand2 gate733( .a(N1588), .b(N2693), .O(N2760) );
buf1 gate734( .a(N2540), .O(N2761) );
buf1 gate735( .a(N2540), .O(N2766) );

  xor2  gate1830(.a(N2695), .b(N2443), .O(gate736inter0));
  nand2 gate1831(.a(gate736inter0), .b(s_80), .O(gate736inter1));
  and2  gate1832(.a(N2695), .b(N2443), .O(gate736inter2));
  inv1  gate1833(.a(s_80), .O(gate736inter3));
  inv1  gate1834(.a(s_81), .O(gate736inter4));
  nand2 gate1835(.a(gate736inter4), .b(gate736inter3), .O(gate736inter5));
  nor2  gate1836(.a(gate736inter5), .b(gate736inter2), .O(gate736inter6));
  inv1  gate1837(.a(N2443), .O(gate736inter7));
  inv1  gate1838(.a(N2695), .O(gate736inter8));
  nand2 gate1839(.a(gate736inter8), .b(gate736inter7), .O(gate736inter9));
  nand2 gate1840(.a(s_81), .b(gate736inter3), .O(gate736inter10));
  nor2  gate1841(.a(gate736inter10), .b(gate736inter9), .O(gate736inter11));
  nor2  gate1842(.a(gate736inter11), .b(gate736inter6), .O(gate736inter12));
  nand2 gate1843(.a(gate736inter12), .b(gate736inter1), .O(N2771));
nand2 gate737( .a(N2440), .b(N2696), .O(N2772) );
nand2 gate738( .a(N2449), .b(N2697), .O(N2773) );

  xor2  gate1494(.a(N2698), .b(N2446), .O(gate739inter0));
  nand2 gate1495(.a(gate739inter0), .b(s_32), .O(gate739inter1));
  and2  gate1496(.a(N2698), .b(N2446), .O(gate739inter2));
  inv1  gate1497(.a(s_32), .O(gate739inter3));
  inv1  gate1498(.a(s_33), .O(gate739inter4));
  nand2 gate1499(.a(gate739inter4), .b(gate739inter3), .O(gate739inter5));
  nor2  gate1500(.a(gate739inter5), .b(gate739inter2), .O(gate739inter6));
  inv1  gate1501(.a(N2446), .O(gate739inter7));
  inv1  gate1502(.a(N2698), .O(gate739inter8));
  nand2 gate1503(.a(gate739inter8), .b(gate739inter7), .O(gate739inter9));
  nand2 gate1504(.a(s_33), .b(gate739inter3), .O(gate739inter10));
  nor2  gate1505(.a(gate739inter10), .b(gate739inter9), .O(gate739inter11));
  nor2  gate1506(.a(gate739inter11), .b(gate739inter6), .O(gate739inter12));
  nand2 gate1507(.a(gate739inter12), .b(gate739inter1), .O(N2774));
nand2 gate740( .a(N2460), .b(N2699), .O(N2775) );
nand2 gate741( .a(N2457), .b(N2700), .O(N2776) );
nand2 gate742( .a(N2466), .b(N2701), .O(N2777) );
nand2 gate743( .a(N2463), .b(N2702), .O(N2778) );
nand2 gate744( .a(N2490), .b(N2707), .O(N2781) );

  xor2  gate1452(.a(N2708), .b(N2487), .O(gate745inter0));
  nand2 gate1453(.a(gate745inter0), .b(s_26), .O(gate745inter1));
  and2  gate1454(.a(N2708), .b(N2487), .O(gate745inter2));
  inv1  gate1455(.a(s_26), .O(gate745inter3));
  inv1  gate1456(.a(s_27), .O(gate745inter4));
  nand2 gate1457(.a(gate745inter4), .b(gate745inter3), .O(gate745inter5));
  nor2  gate1458(.a(gate745inter5), .b(gate745inter2), .O(gate745inter6));
  inv1  gate1459(.a(N2487), .O(gate745inter7));
  inv1  gate1460(.a(N2708), .O(gate745inter8));
  nand2 gate1461(.a(gate745inter8), .b(gate745inter7), .O(gate745inter9));
  nand2 gate1462(.a(s_27), .b(gate745inter3), .O(gate745inter10));
  nor2  gate1463(.a(gate745inter10), .b(gate745inter9), .O(gate745inter11));
  nor2  gate1464(.a(gate745inter11), .b(gate745inter6), .O(gate745inter12));
  nand2 gate1465(.a(gate745inter12), .b(gate745inter1), .O(N2782));
or2 gate746( .a(N2709), .b(N2534), .O(N2783) );
or2 gate747( .a(N2710), .b(N2531), .O(N2784) );
and2 gate748( .a(N1856), .b(N2638), .O(N2789) );
and2 gate749( .a(N1863), .b(N2638), .O(N2790) );
and2 gate750( .a(N1870), .b(N2638), .O(N2791) );
and2 gate751( .a(N1875), .b(N2638), .O(N2792) );
inv1 gate752( .a(N2613), .O(N2793) );

  xor2  gate1438(.a(N2618), .b(N2719), .O(gate753inter0));
  nand2 gate1439(.a(gate753inter0), .b(s_24), .O(gate753inter1));
  and2  gate1440(.a(N2618), .b(N2719), .O(gate753inter2));
  inv1  gate1441(.a(s_24), .O(gate753inter3));
  inv1  gate1442(.a(s_25), .O(gate753inter4));
  nand2 gate1443(.a(gate753inter4), .b(gate753inter3), .O(gate753inter5));
  nor2  gate1444(.a(gate753inter5), .b(gate753inter2), .O(gate753inter6));
  inv1  gate1445(.a(N2719), .O(gate753inter7));
  inv1  gate1446(.a(N2618), .O(gate753inter8));
  nand2 gate1447(.a(gate753inter8), .b(gate753inter7), .O(gate753inter9));
  nand2 gate1448(.a(s_25), .b(gate753inter3), .O(gate753inter10));
  nor2  gate1449(.a(gate753inter10), .b(gate753inter9), .O(gate753inter11));
  nor2  gate1450(.a(gate753inter11), .b(gate753inter6), .O(gate753inter12));
  nand2 gate1451(.a(gate753inter12), .b(gate753inter1), .O(N2796));

  xor2  gate1760(.a(N2720), .b(N2619), .O(gate754inter0));
  nand2 gate1761(.a(gate754inter0), .b(s_70), .O(gate754inter1));
  and2  gate1762(.a(N2720), .b(N2619), .O(gate754inter2));
  inv1  gate1763(.a(s_70), .O(gate754inter3));
  inv1  gate1764(.a(s_71), .O(gate754inter4));
  nand2 gate1765(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate1766(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate1767(.a(N2619), .O(gate754inter7));
  inv1  gate1768(.a(N2720), .O(gate754inter8));
  nand2 gate1769(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate1770(.a(s_71), .b(gate754inter3), .O(gate754inter10));
  nor2  gate1771(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate1772(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate1773(.a(gate754inter12), .b(gate754inter1), .O(N2800));
inv1 gate755( .a(N2624), .O(N2803) );

  xor2  gate1816(.a(N2629), .b(N2726), .O(gate756inter0));
  nand2 gate1817(.a(gate756inter0), .b(s_78), .O(gate756inter1));
  and2  gate1818(.a(N2629), .b(N2726), .O(gate756inter2));
  inv1  gate1819(.a(s_78), .O(gate756inter3));
  inv1  gate1820(.a(s_79), .O(gate756inter4));
  nand2 gate1821(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate1822(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate1823(.a(N2726), .O(gate756inter7));
  inv1  gate1824(.a(N2629), .O(gate756inter8));
  nand2 gate1825(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate1826(.a(s_79), .b(gate756inter3), .O(gate756inter10));
  nor2  gate1827(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate1828(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate1829(.a(gate756inter12), .b(gate756inter1), .O(N2806));
and2 gate757( .a(N1856), .b(N2646), .O(N2809) );
and2 gate758( .a(N1863), .b(N2646), .O(N2810) );
and2 gate759( .a(N1870), .b(N2646), .O(N2811) );
and2 gate760( .a(N1875), .b(N2646), .O(N2812) );
and2 gate761( .a(N2743), .b(N14), .O(N2817) );
buf1 gate762( .a(N2603), .O(N2820) );
nand2 gate763( .a(N2747), .b(N2664), .O(N2826) );
and2 gate764( .a(N2748), .b(N2749), .O(N2829) );
and2 gate765( .a(N2750), .b(N2751), .O(N2830) );
buf1 gate766( .a(N2659), .O(N2831) );
inv1 gate767( .a(N2687), .O(N2837) );
inv1 gate768( .a(N2690), .O(N2838) );
and3 gate769( .a(N2421), .b(N2417), .c(N2687), .O(N2839) );
and3 gate770( .a(N2684), .b(N2681), .c(N2690), .O(N2840) );
nand2 gate771( .a(N2760), .b(N2694), .O(N2841) );
buf1 gate772( .a(N2603), .O(N2844) );
buf1 gate773( .a(N2603), .O(N2854) );
buf1 gate774( .a(N2659), .O(N2859) );
buf1 gate775( .a(N2659), .O(N2869) );
nand2 gate776( .a(N2773), .b(N2774), .O(N2874) );

  xor2  gate2040(.a(N2772), .b(N2771), .O(gate777inter0));
  nand2 gate2041(.a(gate777inter0), .b(s_110), .O(gate777inter1));
  and2  gate2042(.a(N2772), .b(N2771), .O(gate777inter2));
  inv1  gate2043(.a(s_110), .O(gate777inter3));
  inv1  gate2044(.a(s_111), .O(gate777inter4));
  nand2 gate2045(.a(gate777inter4), .b(gate777inter3), .O(gate777inter5));
  nor2  gate2046(.a(gate777inter5), .b(gate777inter2), .O(gate777inter6));
  inv1  gate2047(.a(N2771), .O(gate777inter7));
  inv1  gate2048(.a(N2772), .O(gate777inter8));
  nand2 gate2049(.a(gate777inter8), .b(gate777inter7), .O(gate777inter9));
  nand2 gate2050(.a(s_111), .b(gate777inter3), .O(gate777inter10));
  nor2  gate2051(.a(gate777inter10), .b(gate777inter9), .O(gate777inter11));
  nor2  gate2052(.a(gate777inter11), .b(gate777inter6), .O(gate777inter12));
  nand2 gate2053(.a(gate777inter12), .b(gate777inter1), .O(N2877));
inv1 gate778( .a(N2703), .O(N2880) );
nand2 gate779( .a(N2703), .b(N2706), .O(N2881) );
nand2 gate780( .a(N2777), .b(N2778), .O(N2882) );
nand2 gate781( .a(N2775), .b(N2776), .O(N2885) );
nand2 gate782( .a(N2781), .b(N2782), .O(N2888) );

  xor2  gate1326(.a(N2784), .b(N2783), .O(gate783inter0));
  nand2 gate1327(.a(gate783inter0), .b(s_8), .O(gate783inter1));
  and2  gate1328(.a(N2784), .b(N2783), .O(gate783inter2));
  inv1  gate1329(.a(s_8), .O(gate783inter3));
  inv1  gate1330(.a(s_9), .O(gate783inter4));
  nand2 gate1331(.a(gate783inter4), .b(gate783inter3), .O(gate783inter5));
  nor2  gate1332(.a(gate783inter5), .b(gate783inter2), .O(gate783inter6));
  inv1  gate1333(.a(N2783), .O(gate783inter7));
  inv1  gate1334(.a(N2784), .O(gate783inter8));
  nand2 gate1335(.a(gate783inter8), .b(gate783inter7), .O(gate783inter9));
  nand2 gate1336(.a(s_9), .b(gate783inter3), .O(gate783inter10));
  nor2  gate1337(.a(gate783inter10), .b(gate783inter9), .O(gate783inter11));
  nor2  gate1338(.a(gate783inter11), .b(gate783inter6), .O(gate783inter12));
  nand2 gate1339(.a(gate783inter12), .b(gate783inter1), .O(N2891));
and2 gate784( .a(N2607), .b(N2729), .O(N2894) );
and2 gate785( .a(N2608), .b(N2729), .O(N2895) );
and2 gate786( .a(N2609), .b(N2729), .O(N2896) );
and2 gate787( .a(N2610), .b(N2729), .O(N2897) );
or2 gate788( .a(N2789), .b(N2611), .O(N2898) );
or2 gate789( .a(N2790), .b(N2612), .O(N2899) );
and2 gate790( .a(N2791), .b(N1037), .O(N2900) );
and2 gate791( .a(N2792), .b(N1037), .O(N2901) );
or2 gate792( .a(N2809), .b(N2631), .O(N2914) );
or2 gate793( .a(N2810), .b(N2632), .O(N2915) );
and2 gate794( .a(N2811), .b(N1070), .O(N2916) );
and2 gate795( .a(N2812), .b(N1070), .O(N2917) );
and2 gate796( .a(N2633), .b(N2738), .O(N2918) );
and2 gate797( .a(N2634), .b(N2738), .O(N2919) );
and2 gate798( .a(N2635), .b(N2738), .O(N2920) );
and2 gate799( .a(N2636), .b(N2738), .O(N2921) );
buf1 gate800( .a(N2817), .O(N2925) );
and3 gate801( .a(N2829), .b(N2830), .c(N1302), .O(N2931) );
and3 gate802( .a(N2681), .b(N2421), .c(N2837), .O(N2938) );
and3 gate803( .a(N2417), .b(N2684), .c(N2838), .O(N2939) );
nand2 gate804( .a(N2469), .b(N2880), .O(N2963) );
inv1 gate805( .a(N2841), .O(N2970) );
inv1 gate806( .a(N2826), .O(N2971) );
inv1 gate807( .a(N2894), .O(N2972) );
inv1 gate808( .a(N2895), .O(N2975) );
inv1 gate809( .a(N2896), .O(N2978) );
inv1 gate810( .a(N2897), .O(N2981) );
and2 gate811( .a(N2898), .b(N1037), .O(N2984) );
and2 gate812( .a(N2899), .b(N1037), .O(N2985) );
inv1 gate813( .a(N2900), .O(N2986) );
inv1 gate814( .a(N2901), .O(N2989) );
inv1 gate815( .a(N2796), .O(N2992) );
buf1 gate816( .a(N2800), .O(N2995) );
buf1 gate817( .a(N2800), .O(N2998) );
buf1 gate818( .a(N2806), .O(N3001) );
buf1 gate819( .a(N2806), .O(N3004) );
and2 gate820( .a(N574), .b(N2820), .O(N3007) );
and2 gate821( .a(N2914), .b(N1070), .O(N3008) );
and2 gate822( .a(N2915), .b(N1070), .O(N3009) );
inv1 gate823( .a(N2916), .O(N3010) );
inv1 gate824( .a(N2917), .O(N3013) );
inv1 gate825( .a(N2918), .O(N3016) );
inv1 gate826( .a(N2919), .O(N3019) );
inv1 gate827( .a(N2920), .O(N3022) );
inv1 gate828( .a(N2921), .O(N3025) );
inv1 gate829( .a(N2817), .O(N3028) );
and2 gate830( .a(N574), .b(N2831), .O(N3029) );
inv1 gate831( .a(N2820), .O(N3030) );
and2 gate832( .a(N578), .b(N2820), .O(N3035) );
and2 gate833( .a(N655), .b(N2820), .O(N3036) );
and2 gate834( .a(N659), .b(N2820), .O(N3037) );
buf1 gate835( .a(N2931), .O(N3038) );
inv1 gate836( .a(N2831), .O(N3039) );
and2 gate837( .a(N578), .b(N2831), .O(N3044) );
and2 gate838( .a(N655), .b(N2831), .O(N3045) );
and2 gate839( .a(N659), .b(N2831), .O(N3046) );
nor2 gate840( .a(N2938), .b(N2839), .O(N3047) );
nor2 gate841( .a(N2939), .b(N2840), .O(N3048) );
inv1 gate842( .a(N2888), .O(N3049) );
inv1 gate843( .a(N2844), .O(N3050) );
and2 gate844( .a(N663), .b(N2844), .O(N3053) );
and2 gate845( .a(N667), .b(N2844), .O(N3054) );
and2 gate846( .a(N671), .b(N2844), .O(N3055) );
and2 gate847( .a(N675), .b(N2844), .O(N3056) );
and2 gate848( .a(N679), .b(N2854), .O(N3057) );
and2 gate849( .a(N683), .b(N2854), .O(N3058) );
and2 gate850( .a(N687), .b(N2854), .O(N3059) );
and2 gate851( .a(N705), .b(N2854), .O(N3060) );
inv1 gate852( .a(N2859), .O(N3061) );
and2 gate853( .a(N663), .b(N2859), .O(N3064) );
and2 gate854( .a(N667), .b(N2859), .O(N3065) );
and2 gate855( .a(N671), .b(N2859), .O(N3066) );
and2 gate856( .a(N675), .b(N2859), .O(N3067) );
and2 gate857( .a(N679), .b(N2869), .O(N3068) );
and2 gate858( .a(N683), .b(N2869), .O(N3069) );
and2 gate859( .a(N687), .b(N2869), .O(N3070) );
and2 gate860( .a(N705), .b(N2869), .O(N3071) );
inv1 gate861( .a(N2874), .O(N3072) );
inv1 gate862( .a(N2877), .O(N3073) );
inv1 gate863( .a(N2882), .O(N3074) );
inv1 gate864( .a(N2885), .O(N3075) );

  xor2  gate1508(.a(N2963), .b(N2881), .O(gate865inter0));
  nand2 gate1509(.a(gate865inter0), .b(s_34), .O(gate865inter1));
  and2  gate1510(.a(N2963), .b(N2881), .O(gate865inter2));
  inv1  gate1511(.a(s_34), .O(gate865inter3));
  inv1  gate1512(.a(s_35), .O(gate865inter4));
  nand2 gate1513(.a(gate865inter4), .b(gate865inter3), .O(gate865inter5));
  nor2  gate1514(.a(gate865inter5), .b(gate865inter2), .O(gate865inter6));
  inv1  gate1515(.a(N2881), .O(gate865inter7));
  inv1  gate1516(.a(N2963), .O(gate865inter8));
  nand2 gate1517(.a(gate865inter8), .b(gate865inter7), .O(gate865inter9));
  nand2 gate1518(.a(s_35), .b(gate865inter3), .O(gate865inter10));
  nor2  gate1519(.a(gate865inter10), .b(gate865inter9), .O(gate865inter11));
  nor2  gate1520(.a(gate865inter11), .b(gate865inter6), .O(gate865inter12));
  nand2 gate1521(.a(gate865inter12), .b(gate865inter1), .O(N3076));
inv1 gate866( .a(N2931), .O(N3079) );
inv1 gate867( .a(N2984), .O(N3088) );
inv1 gate868( .a(N2985), .O(N3091) );
inv1 gate869( .a(N3008), .O(N3110) );
inv1 gate870( .a(N3009), .O(N3113) );
and2 gate871( .a(N3055), .b(N1190), .O(N3137) );
and2 gate872( .a(N3056), .b(N1190), .O(N3140) );
and2 gate873( .a(N3057), .b(N2761), .O(N3143) );
and2 gate874( .a(N3058), .b(N2761), .O(N3146) );
and2 gate875( .a(N3059), .b(N2761), .O(N3149) );
and2 gate876( .a(N3060), .b(N2761), .O(N3152) );
and2 gate877( .a(N3066), .b(N1195), .O(N3157) );
and2 gate878( .a(N3067), .b(N1195), .O(N3160) );
and2 gate879( .a(N3068), .b(N2766), .O(N3163) );
and2 gate880( .a(N3069), .b(N2766), .O(N3166) );
and2 gate881( .a(N3070), .b(N2766), .O(N3169) );
and2 gate882( .a(N3071), .b(N2766), .O(N3172) );

  xor2  gate1900(.a(N3072), .b(N2877), .O(gate883inter0));
  nand2 gate1901(.a(gate883inter0), .b(s_90), .O(gate883inter1));
  and2  gate1902(.a(N3072), .b(N2877), .O(gate883inter2));
  inv1  gate1903(.a(s_90), .O(gate883inter3));
  inv1  gate1904(.a(s_91), .O(gate883inter4));
  nand2 gate1905(.a(gate883inter4), .b(gate883inter3), .O(gate883inter5));
  nor2  gate1906(.a(gate883inter5), .b(gate883inter2), .O(gate883inter6));
  inv1  gate1907(.a(N2877), .O(gate883inter7));
  inv1  gate1908(.a(N3072), .O(gate883inter8));
  nand2 gate1909(.a(gate883inter8), .b(gate883inter7), .O(gate883inter9));
  nand2 gate1910(.a(s_91), .b(gate883inter3), .O(gate883inter10));
  nor2  gate1911(.a(gate883inter10), .b(gate883inter9), .O(gate883inter11));
  nor2  gate1912(.a(gate883inter11), .b(gate883inter6), .O(gate883inter12));
  nand2 gate1913(.a(gate883inter12), .b(gate883inter1), .O(N3175));

  xor2  gate1984(.a(N3073), .b(N2874), .O(gate884inter0));
  nand2 gate1985(.a(gate884inter0), .b(s_102), .O(gate884inter1));
  and2  gate1986(.a(N3073), .b(N2874), .O(gate884inter2));
  inv1  gate1987(.a(s_102), .O(gate884inter3));
  inv1  gate1988(.a(s_103), .O(gate884inter4));
  nand2 gate1989(.a(gate884inter4), .b(gate884inter3), .O(gate884inter5));
  nor2  gate1990(.a(gate884inter5), .b(gate884inter2), .O(gate884inter6));
  inv1  gate1991(.a(N2874), .O(gate884inter7));
  inv1  gate1992(.a(N3073), .O(gate884inter8));
  nand2 gate1993(.a(gate884inter8), .b(gate884inter7), .O(gate884inter9));
  nand2 gate1994(.a(s_103), .b(gate884inter3), .O(gate884inter10));
  nor2  gate1995(.a(gate884inter10), .b(gate884inter9), .O(gate884inter11));
  nor2  gate1996(.a(gate884inter11), .b(gate884inter6), .O(gate884inter12));
  nand2 gate1997(.a(gate884inter12), .b(gate884inter1), .O(N3176));

  xor2  gate2026(.a(N3074), .b(N2885), .O(gate885inter0));
  nand2 gate2027(.a(gate885inter0), .b(s_108), .O(gate885inter1));
  and2  gate2028(.a(N3074), .b(N2885), .O(gate885inter2));
  inv1  gate2029(.a(s_108), .O(gate885inter3));
  inv1  gate2030(.a(s_109), .O(gate885inter4));
  nand2 gate2031(.a(gate885inter4), .b(gate885inter3), .O(gate885inter5));
  nor2  gate2032(.a(gate885inter5), .b(gate885inter2), .O(gate885inter6));
  inv1  gate2033(.a(N2885), .O(gate885inter7));
  inv1  gate2034(.a(N3074), .O(gate885inter8));
  nand2 gate2035(.a(gate885inter8), .b(gate885inter7), .O(gate885inter9));
  nand2 gate2036(.a(s_109), .b(gate885inter3), .O(gate885inter10));
  nor2  gate2037(.a(gate885inter10), .b(gate885inter9), .O(gate885inter11));
  nor2  gate2038(.a(gate885inter11), .b(gate885inter6), .O(gate885inter12));
  nand2 gate2039(.a(gate885inter12), .b(gate885inter1), .O(N3177));
nand2 gate886( .a(N2882), .b(N3075), .O(N3178) );
nand2 gate887( .a(N3048), .b(N3047), .O(N3180) );
inv1 gate888( .a(N2995), .O(N3187) );
inv1 gate889( .a(N2998), .O(N3188) );
inv1 gate890( .a(N3001), .O(N3189) );
inv1 gate891( .a(N3004), .O(N3190) );
and3 gate892( .a(N2796), .b(N2613), .c(N2995), .O(N3191) );
and3 gate893( .a(N2992), .b(N2793), .c(N2998), .O(N3192) );
and3 gate894( .a(N2624), .b(N2368), .c(N3001), .O(N3193) );
and3 gate895( .a(N2803), .b(N2621), .c(N3004), .O(N3194) );
nand2 gate896( .a(N3076), .b(N2375), .O(N3195) );
inv1 gate897( .a(N3076), .O(N3196) );
and2 gate898( .a(N687), .b(N3030), .O(N3197) );
and2 gate899( .a(N687), .b(N3039), .O(N3208) );
and2 gate900( .a(N705), .b(N3030), .O(N3215) );
and2 gate901( .a(N711), .b(N3030), .O(N3216) );
and2 gate902( .a(N715), .b(N3030), .O(N3217) );
and2 gate903( .a(N705), .b(N3039), .O(N3218) );
and2 gate904( .a(N711), .b(N3039), .O(N3219) );
and2 gate905( .a(N715), .b(N3039), .O(N3220) );
and2 gate906( .a(N719), .b(N3050), .O(N3222) );
and2 gate907( .a(N723), .b(N3050), .O(N3223) );
and2 gate908( .a(N719), .b(N3061), .O(N3230) );
and2 gate909( .a(N723), .b(N3061), .O(N3231) );
nand2 gate910( .a(N3175), .b(N3176), .O(N3238) );
nand2 gate911( .a(N3177), .b(N3178), .O(N3241) );
buf1 gate912( .a(N2981), .O(N3244) );
buf1 gate913( .a(N2978), .O(N3247) );
buf1 gate914( .a(N2975), .O(N3250) );
buf1 gate915( .a(N2972), .O(N3253) );
buf1 gate916( .a(N2989), .O(N3256) );
buf1 gate917( .a(N2986), .O(N3259) );
buf1 gate918( .a(N3025), .O(N3262) );
buf1 gate919( .a(N3022), .O(N3265) );
buf1 gate920( .a(N3019), .O(N3268) );
buf1 gate921( .a(N3016), .O(N3271) );
buf1 gate922( .a(N3013), .O(N3274) );
buf1 gate923( .a(N3010), .O(N3277) );
and3 gate924( .a(N2793), .b(N2796), .c(N3187), .O(N3281) );
and3 gate925( .a(N2613), .b(N2992), .c(N3188), .O(N3282) );
and3 gate926( .a(N2621), .b(N2624), .c(N3189), .O(N3283) );
and3 gate927( .a(N2368), .b(N2803), .c(N3190), .O(N3284) );
nand2 gate928( .a(N2210), .b(N3196), .O(N3286) );
or2 gate929( .a(N3197), .b(N3007), .O(N3288) );

  xor2  gate1774(.a(N3049), .b(N3180), .O(gate930inter0));
  nand2 gate1775(.a(gate930inter0), .b(s_72), .O(gate930inter1));
  and2  gate1776(.a(N3049), .b(N3180), .O(gate930inter2));
  inv1  gate1777(.a(s_72), .O(gate930inter3));
  inv1  gate1778(.a(s_73), .O(gate930inter4));
  nand2 gate1779(.a(gate930inter4), .b(gate930inter3), .O(gate930inter5));
  nor2  gate1780(.a(gate930inter5), .b(gate930inter2), .O(gate930inter6));
  inv1  gate1781(.a(N3180), .O(gate930inter7));
  inv1  gate1782(.a(N3049), .O(gate930inter8));
  nand2 gate1783(.a(gate930inter8), .b(gate930inter7), .O(gate930inter9));
  nand2 gate1784(.a(s_73), .b(gate930inter3), .O(gate930inter10));
  nor2  gate1785(.a(gate930inter10), .b(gate930inter9), .O(gate930inter11));
  nor2  gate1786(.a(gate930inter11), .b(gate930inter6), .O(gate930inter12));
  nand2 gate1787(.a(gate930inter12), .b(gate930inter1), .O(N3289));
and2 gate931( .a(N3152), .b(N2981), .O(N3291) );
and2 gate932( .a(N3149), .b(N2978), .O(N3293) );
and2 gate933( .a(N3146), .b(N2975), .O(N3295) );
and2 gate934( .a(N2972), .b(N3143), .O(N3296) );
and2 gate935( .a(N3140), .b(N2989), .O(N3299) );
and2 gate936( .a(N3137), .b(N2986), .O(N3301) );
or2 gate937( .a(N3208), .b(N3029), .O(N3302) );
and2 gate938( .a(N3172), .b(N3025), .O(N3304) );
and2 gate939( .a(N3169), .b(N3022), .O(N3306) );
and2 gate940( .a(N3166), .b(N3019), .O(N3308) );
and2 gate941( .a(N3016), .b(N3163), .O(N3309) );
and2 gate942( .a(N3160), .b(N3013), .O(N3312) );
and2 gate943( .a(N3157), .b(N3010), .O(N3314) );
or2 gate944( .a(N3215), .b(N3035), .O(N3315) );
or2 gate945( .a(N3216), .b(N3036), .O(N3318) );
or2 gate946( .a(N3217), .b(N3037), .O(N3321) );
or2 gate947( .a(N3218), .b(N3044), .O(N3324) );
or2 gate948( .a(N3219), .b(N3045), .O(N3327) );
or2 gate949( .a(N3220), .b(N3046), .O(N3330) );
inv1 gate950( .a(N3180), .O(N3333) );
or2 gate951( .a(N3222), .b(N3053), .O(N3334) );
or2 gate952( .a(N3223), .b(N3054), .O(N3335) );
or2 gate953( .a(N3230), .b(N3064), .O(N3336) );
or2 gate954( .a(N3231), .b(N3065), .O(N3337) );
buf1 gate955( .a(N3152), .O(N3340) );
buf1 gate956( .a(N3149), .O(N3344) );
buf1 gate957( .a(N3146), .O(N3348) );
buf1 gate958( .a(N3143), .O(N3352) );
buf1 gate959( .a(N3140), .O(N3356) );
buf1 gate960( .a(N3137), .O(N3360) );
buf1 gate961( .a(N3091), .O(N3364) );
buf1 gate962( .a(N3088), .O(N3367) );
buf1 gate963( .a(N3172), .O(N3370) );
buf1 gate964( .a(N3169), .O(N3374) );
buf1 gate965( .a(N3166), .O(N3378) );
buf1 gate966( .a(N3163), .O(N3382) );
buf1 gate967( .a(N3160), .O(N3386) );
buf1 gate968( .a(N3157), .O(N3390) );
buf1 gate969( .a(N3113), .O(N3394) );
buf1 gate970( .a(N3110), .O(N3397) );
nand2 gate971( .a(N3195), .b(N3286), .O(N3400) );
nor2 gate972( .a(N3281), .b(N3191), .O(N3401) );
nor2 gate973( .a(N3282), .b(N3192), .O(N3402) );
nor2 gate974( .a(N3283), .b(N3193), .O(N3403) );
nor2 gate975( .a(N3284), .b(N3194), .O(N3404) );
inv1 gate976( .a(N3238), .O(N3405) );
inv1 gate977( .a(N3241), .O(N3406) );
and2 gate978( .a(N3288), .b(N1836), .O(N3409) );
nand2 gate979( .a(N2888), .b(N3333), .O(N3410) );
inv1 gate980( .a(N3244), .O(N3412) );
inv1 gate981( .a(N3247), .O(N3414) );
inv1 gate982( .a(N3250), .O(N3416) );
inv1 gate983( .a(N3253), .O(N3418) );
inv1 gate984( .a(N3256), .O(N3420) );
inv1 gate985( .a(N3259), .O(N3422) );
and2 gate986( .a(N3302), .b(N1836), .O(N3428) );
inv1 gate987( .a(N3262), .O(N3430) );
inv1 gate988( .a(N3265), .O(N3432) );
inv1 gate989( .a(N3268), .O(N3434) );
inv1 gate990( .a(N3271), .O(N3436) );
inv1 gate991( .a(N3274), .O(N3438) );
inv1 gate992( .a(N3277), .O(N3440) );
and2 gate993( .a(N3334), .b(N1190), .O(N3450) );
and2 gate994( .a(N3335), .b(N1190), .O(N3453) );
and2 gate995( .a(N3336), .b(N1195), .O(N3456) );
and2 gate996( .a(N3337), .b(N1195), .O(N3459) );
and2 gate997( .a(N3400), .b(N533), .O(N3478) );
and2 gate998( .a(N3318), .b(N2128), .O(N3479) );
and2 gate999( .a(N3315), .b(N1841), .O(N3480) );
nand2 gate1000( .a(N3410), .b(N3289), .O(N3481) );
inv1 gate1001( .a(N3340), .O(N3482) );
nand2 gate1002( .a(N3340), .b(N3412), .O(N3483) );
inv1 gate1003( .a(N3344), .O(N3484) );
nand2 gate1004( .a(N3344), .b(N3414), .O(N3485) );
inv1 gate1005( .a(N3348), .O(N3486) );
nand2 gate1006( .a(N3348), .b(N3416), .O(N3487) );
inv1 gate1007( .a(N3352), .O(N3488) );
nand2 gate1008( .a(N3352), .b(N3418), .O(N3489) );
inv1 gate1009( .a(N3356), .O(N3490) );
nand2 gate1010( .a(N3356), .b(N3420), .O(N3491) );
inv1 gate1011( .a(N3360), .O(N3492) );
nand2 gate1012( .a(N3360), .b(N3422), .O(N3493) );
inv1 gate1013( .a(N3364), .O(N3494) );
inv1 gate1014( .a(N3367), .O(N3496) );
and2 gate1015( .a(N3321), .b(N2135), .O(N3498) );
and2 gate1016( .a(N3327), .b(N2128), .O(N3499) );
and2 gate1017( .a(N3324), .b(N1841), .O(N3500) );
inv1 gate1018( .a(N3370), .O(N3501) );
nand2 gate1019( .a(N3370), .b(N3430), .O(N3502) );
inv1 gate1020( .a(N3374), .O(N3503) );
nand2 gate1021( .a(N3374), .b(N3432), .O(N3504) );
inv1 gate1022( .a(N3378), .O(N3505) );
nand2 gate1023( .a(N3378), .b(N3434), .O(N3506) );
inv1 gate1024( .a(N3382), .O(N3507) );
nand2 gate1025( .a(N3382), .b(N3436), .O(N3508) );
inv1 gate1026( .a(N3386), .O(N3509) );
nand2 gate1027( .a(N3386), .b(N3438), .O(N3510) );
inv1 gate1028( .a(N3390), .O(N3511) );
nand2 gate1029( .a(N3390), .b(N3440), .O(N3512) );
inv1 gate1030( .a(N3394), .O(N3513) );
inv1 gate1031( .a(N3397), .O(N3515) );
and2 gate1032( .a(N3330), .b(N2135), .O(N3517) );
nand2 gate1033( .a(N3402), .b(N3401), .O(N3522) );
nand2 gate1034( .a(N3404), .b(N3403), .O(N3525) );
buf1 gate1035( .a(N3318), .O(N3528) );
buf1 gate1036( .a(N3315), .O(N3531) );
buf1 gate1037( .a(N3321), .O(N3534) );
buf1 gate1038( .a(N3327), .O(N3537) );
buf1 gate1039( .a(N3324), .O(N3540) );
buf1 gate1040( .a(N3330), .O(N3543) );
or2 gate1041( .a(N3478), .b(N1813), .O(N3546) );
inv1 gate1042( .a(N3481), .O(N3551) );
nand2 gate1043( .a(N3244), .b(N3482), .O(N3552) );
nand2 gate1044( .a(N3247), .b(N3484), .O(N3553) );
nand2 gate1045( .a(N3250), .b(N3486), .O(N3554) );
nand2 gate1046( .a(N3253), .b(N3488), .O(N3555) );
nand2 gate1047( .a(N3256), .b(N3490), .O(N3556) );
nand2 gate1048( .a(N3259), .b(N3492), .O(N3557) );
and2 gate1049( .a(N3453), .b(N3091), .O(N3558) );
and2 gate1050( .a(N3450), .b(N3088), .O(N3559) );

  xor2  gate1676(.a(N3501), .b(N3262), .O(gate1051inter0));
  nand2 gate1677(.a(gate1051inter0), .b(s_58), .O(gate1051inter1));
  and2  gate1678(.a(N3501), .b(N3262), .O(gate1051inter2));
  inv1  gate1679(.a(s_58), .O(gate1051inter3));
  inv1  gate1680(.a(s_59), .O(gate1051inter4));
  nand2 gate1681(.a(gate1051inter4), .b(gate1051inter3), .O(gate1051inter5));
  nor2  gate1682(.a(gate1051inter5), .b(gate1051inter2), .O(gate1051inter6));
  inv1  gate1683(.a(N3262), .O(gate1051inter7));
  inv1  gate1684(.a(N3501), .O(gate1051inter8));
  nand2 gate1685(.a(gate1051inter8), .b(gate1051inter7), .O(gate1051inter9));
  nand2 gate1686(.a(s_59), .b(gate1051inter3), .O(gate1051inter10));
  nor2  gate1687(.a(gate1051inter10), .b(gate1051inter9), .O(gate1051inter11));
  nor2  gate1688(.a(gate1051inter11), .b(gate1051inter6), .O(gate1051inter12));
  nand2 gate1689(.a(gate1051inter12), .b(gate1051inter1), .O(N3563));
nand2 gate1052( .a(N3265), .b(N3503), .O(N3564) );
nand2 gate1053( .a(N3268), .b(N3505), .O(N3565) );
nand2 gate1054( .a(N3271), .b(N3507), .O(N3566) );
nand2 gate1055( .a(N3274), .b(N3509), .O(N3567) );

  xor2  gate1704(.a(N3511), .b(N3277), .O(gate1056inter0));
  nand2 gate1705(.a(gate1056inter0), .b(s_62), .O(gate1056inter1));
  and2  gate1706(.a(N3511), .b(N3277), .O(gate1056inter2));
  inv1  gate1707(.a(s_62), .O(gate1056inter3));
  inv1  gate1708(.a(s_63), .O(gate1056inter4));
  nand2 gate1709(.a(gate1056inter4), .b(gate1056inter3), .O(gate1056inter5));
  nor2  gate1710(.a(gate1056inter5), .b(gate1056inter2), .O(gate1056inter6));
  inv1  gate1711(.a(N3277), .O(gate1056inter7));
  inv1  gate1712(.a(N3511), .O(gate1056inter8));
  nand2 gate1713(.a(gate1056inter8), .b(gate1056inter7), .O(gate1056inter9));
  nand2 gate1714(.a(s_63), .b(gate1056inter3), .O(gate1056inter10));
  nor2  gate1715(.a(gate1056inter10), .b(gate1056inter9), .O(gate1056inter11));
  nor2  gate1716(.a(gate1056inter11), .b(gate1056inter6), .O(gate1056inter12));
  nand2 gate1717(.a(gate1056inter12), .b(gate1056inter1), .O(N3568));
and2 gate1057( .a(N3459), .b(N3113), .O(N3569) );
and2 gate1058( .a(N3456), .b(N3110), .O(N3570) );
buf1 gate1059( .a(N3453), .O(N3576) );
buf1 gate1060( .a(N3450), .O(N3579) );
buf1 gate1061( .a(N3459), .O(N3585) );
buf1 gate1062( .a(N3456), .O(N3588) );
inv1 gate1063( .a(N3522), .O(N3592) );
nand2 gate1064( .a(N3522), .b(N3405), .O(N3593) );
inv1 gate1065( .a(N3525), .O(N3594) );
nand2 gate1066( .a(N3525), .b(N3406), .O(N3595) );
inv1 gate1067( .a(N3528), .O(N3596) );
nand2 gate1068( .a(N3528), .b(N2630), .O(N3597) );

  xor2  gate1536(.a(N2376), .b(N3531), .O(gate1069inter0));
  nand2 gate1537(.a(gate1069inter0), .b(s_38), .O(gate1069inter1));
  and2  gate1538(.a(N2376), .b(N3531), .O(gate1069inter2));
  inv1  gate1539(.a(s_38), .O(gate1069inter3));
  inv1  gate1540(.a(s_39), .O(gate1069inter4));
  nand2 gate1541(.a(gate1069inter4), .b(gate1069inter3), .O(gate1069inter5));
  nor2  gate1542(.a(gate1069inter5), .b(gate1069inter2), .O(gate1069inter6));
  inv1  gate1543(.a(N3531), .O(gate1069inter7));
  inv1  gate1544(.a(N2376), .O(gate1069inter8));
  nand2 gate1545(.a(gate1069inter8), .b(gate1069inter7), .O(gate1069inter9));
  nand2 gate1546(.a(s_39), .b(gate1069inter3), .O(gate1069inter10));
  nor2  gate1547(.a(gate1069inter10), .b(gate1069inter9), .O(gate1069inter11));
  nor2  gate1548(.a(gate1069inter11), .b(gate1069inter6), .O(gate1069inter12));
  nand2 gate1549(.a(gate1069inter12), .b(gate1069inter1), .O(N3598));
inv1 gate1070( .a(N3531), .O(N3599) );
and2 gate1071( .a(N3551), .b(N800), .O(N3600) );
nand2 gate1072( .a(N3552), .b(N3483), .O(N3603) );
nand2 gate1073( .a(N3553), .b(N3485), .O(N3608) );
nand2 gate1074( .a(N3554), .b(N3487), .O(N3612) );
nand2 gate1075( .a(N3555), .b(N3489), .O(N3615) );
nand2 gate1076( .a(N3556), .b(N3491), .O(N3616) );
nand2 gate1077( .a(N3557), .b(N3493), .O(N3622) );
inv1 gate1078( .a(N3534), .O(N3629) );

  xor2  gate1606(.a(N2645), .b(N3534), .O(gate1079inter0));
  nand2 gate1607(.a(gate1079inter0), .b(s_48), .O(gate1079inter1));
  and2  gate1608(.a(N2645), .b(N3534), .O(gate1079inter2));
  inv1  gate1609(.a(s_48), .O(gate1079inter3));
  inv1  gate1610(.a(s_49), .O(gate1079inter4));
  nand2 gate1611(.a(gate1079inter4), .b(gate1079inter3), .O(gate1079inter5));
  nor2  gate1612(.a(gate1079inter5), .b(gate1079inter2), .O(gate1079inter6));
  inv1  gate1613(.a(N3534), .O(gate1079inter7));
  inv1  gate1614(.a(N2645), .O(gate1079inter8));
  nand2 gate1615(.a(gate1079inter8), .b(gate1079inter7), .O(gate1079inter9));
  nand2 gate1616(.a(s_49), .b(gate1079inter3), .O(gate1079inter10));
  nor2  gate1617(.a(gate1079inter10), .b(gate1079inter9), .O(gate1079inter11));
  nor2  gate1618(.a(gate1079inter11), .b(gate1079inter6), .O(gate1079inter12));
  nand2 gate1619(.a(gate1079inter12), .b(gate1079inter1), .O(N3630));
inv1 gate1080( .a(N3537), .O(N3631) );

  xor2  gate1312(.a(N2655), .b(N3537), .O(gate1081inter0));
  nand2 gate1313(.a(gate1081inter0), .b(s_6), .O(gate1081inter1));
  and2  gate1314(.a(N2655), .b(N3537), .O(gate1081inter2));
  inv1  gate1315(.a(s_6), .O(gate1081inter3));
  inv1  gate1316(.a(s_7), .O(gate1081inter4));
  nand2 gate1317(.a(gate1081inter4), .b(gate1081inter3), .O(gate1081inter5));
  nor2  gate1318(.a(gate1081inter5), .b(gate1081inter2), .O(gate1081inter6));
  inv1  gate1319(.a(N3537), .O(gate1081inter7));
  inv1  gate1320(.a(N2655), .O(gate1081inter8));
  nand2 gate1321(.a(gate1081inter8), .b(gate1081inter7), .O(gate1081inter9));
  nand2 gate1322(.a(s_7), .b(gate1081inter3), .O(gate1081inter10));
  nor2  gate1323(.a(gate1081inter10), .b(gate1081inter9), .O(gate1081inter11));
  nor2  gate1324(.a(gate1081inter11), .b(gate1081inter6), .O(gate1081inter12));
  nand2 gate1325(.a(gate1081inter12), .b(gate1081inter1), .O(N3632));
nand2 gate1082( .a(N3540), .b(N2403), .O(N3633) );
inv1 gate1083( .a(N3540), .O(N3634) );
nand2 gate1084( .a(N3563), .b(N3502), .O(N3635) );
nand2 gate1085( .a(N3564), .b(N3504), .O(N3640) );
nand2 gate1086( .a(N3565), .b(N3506), .O(N3644) );
nand2 gate1087( .a(N3566), .b(N3508), .O(N3647) );
nand2 gate1088( .a(N3567), .b(N3510), .O(N3648) );
nand2 gate1089( .a(N3568), .b(N3512), .O(N3654) );
inv1 gate1090( .a(N3543), .O(N3661) );
nand2 gate1091( .a(N3543), .b(N2656), .O(N3662) );
nand2 gate1092( .a(N3238), .b(N3592), .O(N3667) );
nand2 gate1093( .a(N3241), .b(N3594), .O(N3668) );
nand2 gate1094( .a(N2472), .b(N3596), .O(N3669) );
nand2 gate1095( .a(N2213), .b(N3599), .O(N3670) );
buf1 gate1096( .a(N3600), .O(N3671) );
inv1 gate1097( .a(N3576), .O(N3691) );
nand2 gate1098( .a(N3576), .b(N3494), .O(N3692) );
inv1 gate1099( .a(N3579), .O(N3693) );
nand2 gate1100( .a(N3579), .b(N3496), .O(N3694) );
nand2 gate1101( .a(N2475), .b(N3629), .O(N3695) );
nand2 gate1102( .a(N2478), .b(N3631), .O(N3696) );
nand2 gate1103( .a(N2216), .b(N3634), .O(N3697) );
inv1 gate1104( .a(N3585), .O(N3716) );

  xor2  gate1690(.a(N3513), .b(N3585), .O(gate1105inter0));
  nand2 gate1691(.a(gate1105inter0), .b(s_60), .O(gate1105inter1));
  and2  gate1692(.a(N3513), .b(N3585), .O(gate1105inter2));
  inv1  gate1693(.a(s_60), .O(gate1105inter3));
  inv1  gate1694(.a(s_61), .O(gate1105inter4));
  nand2 gate1695(.a(gate1105inter4), .b(gate1105inter3), .O(gate1105inter5));
  nor2  gate1696(.a(gate1105inter5), .b(gate1105inter2), .O(gate1105inter6));
  inv1  gate1697(.a(N3585), .O(gate1105inter7));
  inv1  gate1698(.a(N3513), .O(gate1105inter8));
  nand2 gate1699(.a(gate1105inter8), .b(gate1105inter7), .O(gate1105inter9));
  nand2 gate1700(.a(s_61), .b(gate1105inter3), .O(gate1105inter10));
  nor2  gate1701(.a(gate1105inter10), .b(gate1105inter9), .O(gate1105inter11));
  nor2  gate1702(.a(gate1105inter11), .b(gate1105inter6), .O(gate1105inter12));
  nand2 gate1703(.a(gate1105inter12), .b(gate1105inter1), .O(N3717));
inv1 gate1106( .a(N3588), .O(N3718) );
nand2 gate1107( .a(N3588), .b(N3515), .O(N3719) );
nand2 gate1108( .a(N2481), .b(N3661), .O(N3720) );
nand2 gate1109( .a(N3667), .b(N3593), .O(N3721) );
nand2 gate1110( .a(N3668), .b(N3595), .O(N3722) );
nand2 gate1111( .a(N3669), .b(N3597), .O(N3723) );
nand2 gate1112( .a(N3670), .b(N3598), .O(N3726) );
inv1 gate1113( .a(N3600), .O(N3727) );
nand2 gate1114( .a(N3364), .b(N3691), .O(N3728) );
nand2 gate1115( .a(N3367), .b(N3693), .O(N3729) );

  xor2  gate1340(.a(N3630), .b(N3695), .O(gate1116inter0));
  nand2 gate1341(.a(gate1116inter0), .b(s_10), .O(gate1116inter1));
  and2  gate1342(.a(N3630), .b(N3695), .O(gate1116inter2));
  inv1  gate1343(.a(s_10), .O(gate1116inter3));
  inv1  gate1344(.a(s_11), .O(gate1116inter4));
  nand2 gate1345(.a(gate1116inter4), .b(gate1116inter3), .O(gate1116inter5));
  nor2  gate1346(.a(gate1116inter5), .b(gate1116inter2), .O(gate1116inter6));
  inv1  gate1347(.a(N3695), .O(gate1116inter7));
  inv1  gate1348(.a(N3630), .O(gate1116inter8));
  nand2 gate1349(.a(gate1116inter8), .b(gate1116inter7), .O(gate1116inter9));
  nand2 gate1350(.a(s_11), .b(gate1116inter3), .O(gate1116inter10));
  nor2  gate1351(.a(gate1116inter10), .b(gate1116inter9), .O(gate1116inter11));
  nor2  gate1352(.a(gate1116inter11), .b(gate1116inter6), .O(gate1116inter12));
  nand2 gate1353(.a(gate1116inter12), .b(gate1116inter1), .O(N3730));
and4 gate1117( .a(N3608), .b(N3615), .c(N3612), .d(N3603), .O(N3731) );
and2 gate1118( .a(N3603), .b(N3293), .O(N3732) );
and3 gate1119( .a(N3608), .b(N3603), .c(N3295), .O(N3733) );
and4 gate1120( .a(N3612), .b(N3603), .c(N3296), .d(N3608), .O(N3734) );
and2 gate1121( .a(N3616), .b(N3301), .O(N3735) );
and3 gate1122( .a(N3622), .b(N3616), .c(N3558), .O(N3736) );
nand2 gate1123( .a(N3696), .b(N3632), .O(N3737) );
nand2 gate1124( .a(N3697), .b(N3633), .O(N3740) );
nand2 gate1125( .a(N3394), .b(N3716), .O(N3741) );

  xor2  gate1788(.a(N3718), .b(N3397), .O(gate1126inter0));
  nand2 gate1789(.a(gate1126inter0), .b(s_74), .O(gate1126inter1));
  and2  gate1790(.a(N3718), .b(N3397), .O(gate1126inter2));
  inv1  gate1791(.a(s_74), .O(gate1126inter3));
  inv1  gate1792(.a(s_75), .O(gate1126inter4));
  nand2 gate1793(.a(gate1126inter4), .b(gate1126inter3), .O(gate1126inter5));
  nor2  gate1794(.a(gate1126inter5), .b(gate1126inter2), .O(gate1126inter6));
  inv1  gate1795(.a(N3397), .O(gate1126inter7));
  inv1  gate1796(.a(N3718), .O(gate1126inter8));
  nand2 gate1797(.a(gate1126inter8), .b(gate1126inter7), .O(gate1126inter9));
  nand2 gate1798(.a(s_75), .b(gate1126inter3), .O(gate1126inter10));
  nor2  gate1799(.a(gate1126inter10), .b(gate1126inter9), .O(gate1126inter11));
  nor2  gate1800(.a(gate1126inter11), .b(gate1126inter6), .O(gate1126inter12));
  nand2 gate1801(.a(gate1126inter12), .b(gate1126inter1), .O(N3742));
nand2 gate1127( .a(N3720), .b(N3662), .O(N3743) );
and4 gate1128( .a(N3640), .b(N3647), .c(N3644), .d(N3635), .O(N3744) );
and2 gate1129( .a(N3635), .b(N3306), .O(N3745) );
and3 gate1130( .a(N3640), .b(N3635), .c(N3308), .O(N3746) );
and4 gate1131( .a(N3644), .b(N3635), .c(N3309), .d(N3640), .O(N3747) );
and2 gate1132( .a(N3648), .b(N3314), .O(N3748) );
and3 gate1133( .a(N3654), .b(N3648), .c(N3569), .O(N3749) );
inv1 gate1134( .a(N3721), .O(N3750) );
and2 gate1135( .a(N3722), .b(N246), .O(N3753) );
nand2 gate1136( .a(N3728), .b(N3692), .O(N3754) );
nand2 gate1137( .a(N3729), .b(N3694), .O(N3758) );
inv1 gate1138( .a(N3731), .O(N3761) );
or4 gate1139( .a(N3291), .b(N3732), .c(N3733), .d(N3734), .O(N3762) );
nand2 gate1140( .a(N3741), .b(N3717), .O(N3767) );

  xor2  gate1634(.a(N3719), .b(N3742), .O(gate1141inter0));
  nand2 gate1635(.a(gate1141inter0), .b(s_52), .O(gate1141inter1));
  and2  gate1636(.a(N3719), .b(N3742), .O(gate1141inter2));
  inv1  gate1637(.a(s_52), .O(gate1141inter3));
  inv1  gate1638(.a(s_53), .O(gate1141inter4));
  nand2 gate1639(.a(gate1141inter4), .b(gate1141inter3), .O(gate1141inter5));
  nor2  gate1640(.a(gate1141inter5), .b(gate1141inter2), .O(gate1141inter6));
  inv1  gate1641(.a(N3742), .O(gate1141inter7));
  inv1  gate1642(.a(N3719), .O(gate1141inter8));
  nand2 gate1643(.a(gate1141inter8), .b(gate1141inter7), .O(gate1141inter9));
  nand2 gate1644(.a(s_53), .b(gate1141inter3), .O(gate1141inter10));
  nor2  gate1645(.a(gate1141inter10), .b(gate1141inter9), .O(gate1141inter11));
  nor2  gate1646(.a(gate1141inter11), .b(gate1141inter6), .O(gate1141inter12));
  nand2 gate1647(.a(gate1141inter12), .b(gate1141inter1), .O(N3771));
inv1 gate1142( .a(N3744), .O(N3774) );
or4 gate1143( .a(N3304), .b(N3745), .c(N3746), .d(N3747), .O(N3775) );
and2 gate1144( .a(N3723), .b(N3480), .O(N3778) );
and3 gate1145( .a(N3726), .b(N3723), .c(N3409), .O(N3779) );
or2 gate1146( .a(N2125), .b(N3753), .O(N3780) );
and2 gate1147( .a(N3750), .b(N800), .O(N3790) );
and2 gate1148( .a(N3737), .b(N3500), .O(N3793) );
and3 gate1149( .a(N3740), .b(N3737), .c(N3428), .O(N3794) );
or3 gate1150( .a(N3479), .b(N3778), .c(N3779), .O(N3802) );
buf1 gate1151( .a(N3780), .O(N3803) );
buf1 gate1152( .a(N3780), .O(N3804) );
inv1 gate1153( .a(N3762), .O(N3805) );
and5 gate1154( .a(N3622), .b(N3730), .c(N3754), .d(N3616), .e(N3758), .O(N3806) );
and4 gate1155( .a(N3754), .b(N3616), .c(N3559), .d(N3622), .O(N3807) );
and5 gate1156( .a(N3758), .b(N3754), .c(N3616), .d(N3498), .e(N3622), .O(N3808) );
buf1 gate1157( .a(N3790), .O(N3809) );
or3 gate1158( .a(N3499), .b(N3793), .c(N3794), .O(N3811) );
inv1 gate1159( .a(N3775), .O(N3812) );
and5 gate1160( .a(N3654), .b(N3743), .c(N3767), .d(N3648), .e(N3771), .O(N3813) );
and4 gate1161( .a(N3767), .b(N3648), .c(N3570), .d(N3654), .O(N3814) );
and5 gate1162( .a(N3771), .b(N3767), .c(N3648), .d(N3517), .e(N3654), .O(N3815) );
or5 gate1163( .a(N3299), .b(N3735), .c(N3736), .d(N3807), .e(N3808), .O(N3816) );
and2 gate1164( .a(N3806), .b(N3802), .O(N3817) );
nand2 gate1165( .a(N3805), .b(N3761), .O(N3818) );
inv1 gate1166( .a(N3790), .O(N3819) );
or5 gate1167( .a(N3312), .b(N3748), .c(N3749), .d(N3814), .e(N3815), .O(N3820) );
and2 gate1168( .a(N3813), .b(N3811), .O(N3821) );

  xor2  gate1858(.a(N3774), .b(N3812), .O(gate1169inter0));
  nand2 gate1859(.a(gate1169inter0), .b(s_84), .O(gate1169inter1));
  and2  gate1860(.a(N3774), .b(N3812), .O(gate1169inter2));
  inv1  gate1861(.a(s_84), .O(gate1169inter3));
  inv1  gate1862(.a(s_85), .O(gate1169inter4));
  nand2 gate1863(.a(gate1169inter4), .b(gate1169inter3), .O(gate1169inter5));
  nor2  gate1864(.a(gate1169inter5), .b(gate1169inter2), .O(gate1169inter6));
  inv1  gate1865(.a(N3812), .O(gate1169inter7));
  inv1  gate1866(.a(N3774), .O(gate1169inter8));
  nand2 gate1867(.a(gate1169inter8), .b(gate1169inter7), .O(gate1169inter9));
  nand2 gate1868(.a(s_85), .b(gate1169inter3), .O(gate1169inter10));
  nor2  gate1869(.a(gate1169inter10), .b(gate1169inter9), .O(gate1169inter11));
  nor2  gate1870(.a(gate1169inter11), .b(gate1169inter6), .O(gate1169inter12));
  nand2 gate1871(.a(gate1169inter12), .b(gate1169inter1), .O(N3822));
or2 gate1170( .a(N3816), .b(N3817), .O(N3823) );
and3 gate1171( .a(N3727), .b(N3819), .c(N2841), .O(N3826) );
or2 gate1172( .a(N3820), .b(N3821), .O(N3827) );
inv1 gate1173( .a(N3823), .O(N3834) );
and2 gate1174( .a(N3818), .b(N3823), .O(N3835) );
inv1 gate1175( .a(N3827), .O(N3836) );
and2 gate1176( .a(N3822), .b(N3827), .O(N3837) );
and2 gate1177( .a(N3762), .b(N3834), .O(N3838) );
and2 gate1178( .a(N3775), .b(N3836), .O(N3839) );
or2 gate1179( .a(N3838), .b(N3835), .O(N3840) );
or2 gate1180( .a(N3839), .b(N3837), .O(N3843) );
buf1 gate1181( .a(N3843), .O(N3851) );

  xor2  gate1746(.a(N3840), .b(N3843), .O(gate1182inter0));
  nand2 gate1747(.a(gate1182inter0), .b(s_68), .O(gate1182inter1));
  and2  gate1748(.a(N3840), .b(N3843), .O(gate1182inter2));
  inv1  gate1749(.a(s_68), .O(gate1182inter3));
  inv1  gate1750(.a(s_69), .O(gate1182inter4));
  nand2 gate1751(.a(gate1182inter4), .b(gate1182inter3), .O(gate1182inter5));
  nor2  gate1752(.a(gate1182inter5), .b(gate1182inter2), .O(gate1182inter6));
  inv1  gate1753(.a(N3843), .O(gate1182inter7));
  inv1  gate1754(.a(N3840), .O(gate1182inter8));
  nand2 gate1755(.a(gate1182inter8), .b(gate1182inter7), .O(gate1182inter9));
  nand2 gate1756(.a(s_69), .b(gate1182inter3), .O(gate1182inter10));
  nor2  gate1757(.a(gate1182inter10), .b(gate1182inter9), .O(gate1182inter11));
  nor2  gate1758(.a(gate1182inter11), .b(gate1182inter6), .O(gate1182inter12));
  nand2 gate1759(.a(gate1182inter12), .b(gate1182inter1), .O(N3852));
and2 gate1183( .a(N3843), .b(N3852), .O(N3857) );
and2 gate1184( .a(N3852), .b(N3840), .O(N3858) );
or2 gate1185( .a(N3857), .b(N3858), .O(N3859) );
inv1 gate1186( .a(N3859), .O(N3864) );
and2 gate1187( .a(N3859), .b(N3864), .O(N3869) );
or2 gate1188( .a(N3869), .b(N3864), .O(N3870) );
inv1 gate1189( .a(N3870), .O(N3875) );
and3 gate1190( .a(N2826), .b(N3028), .c(N3870), .O(N3876) );
and3 gate1191( .a(N3826), .b(N3876), .c(N1591), .O(N3877) );
buf1 gate1192( .a(N3877), .O(N3881) );
inv1 gate1193( .a(N3877), .O(N3882) );
buf1 gate1194( .a(N143_I), .O(N143_O) );
buf1 gate1195( .a(N144_I), .O(N144_O) );
buf1 gate1196( .a(N145_I), .O(N145_O) );
buf1 gate1197( .a(N146_I), .O(N146_O) );
buf1 gate1198( .a(N147_I), .O(N147_O) );
buf1 gate1199( .a(N148_I), .O(N148_O) );
buf1 gate1200( .a(N149_I), .O(N149_O) );
buf1 gate1201( .a(N150_I), .O(N150_O) );
buf1 gate1202( .a(N151_I), .O(N151_O) );
buf1 gate1203( .a(N152_I), .O(N152_O) );
buf1 gate1204( .a(N153_I), .O(N153_O) );
buf1 gate1205( .a(N154_I), .O(N154_O) );
buf1 gate1206( .a(N155_I), .O(N155_O) );
buf1 gate1207( .a(N156_I), .O(N156_O) );
buf1 gate1208( .a(N157_I), .O(N157_O) );
buf1 gate1209( .a(N158_I), .O(N158_O) );
buf1 gate1210( .a(N159_I), .O(N159_O) );
buf1 gate1211( .a(N160_I), .O(N160_O) );
buf1 gate1212( .a(N161_I), .O(N161_O) );
buf1 gate1213( .a(N162_I), .O(N162_O) );
buf1 gate1214( .a(N163_I), .O(N163_O) );
buf1 gate1215( .a(N164_I), .O(N164_O) );
buf1 gate1216( .a(N165_I), .O(N165_O) );
buf1 gate1217( .a(N166_I), .O(N166_O) );
buf1 gate1218( .a(N167_I), .O(N167_O) );
buf1 gate1219( .a(N168_I), .O(N168_O) );
buf1 gate1220( .a(N169_I), .O(N169_O) );
buf1 gate1221( .a(N170_I), .O(N170_O) );
buf1 gate1222( .a(N171_I), .O(N171_O) );
buf1 gate1223( .a(N172_I), .O(N172_O) );
buf1 gate1224( .a(N173_I), .O(N173_O) );
buf1 gate1225( .a(N174_I), .O(N174_O) );
buf1 gate1226( .a(N175_I), .O(N175_O) );
buf1 gate1227( .a(N176_I), .O(N176_O) );
buf1 gate1228( .a(N177_I), .O(N177_O) );
buf1 gate1229( .a(N178_I), .O(N178_O) );
buf1 gate1230( .a(N179_I), .O(N179_O) );
buf1 gate1231( .a(N180_I), .O(N180_O) );
buf1 gate1232( .a(N181_I), .O(N181_O) );
buf1 gate1233( .a(N182_I), .O(N182_O) );
buf1 gate1234( .a(N183_I), .O(N183_O) );
buf1 gate1235( .a(N184_I), .O(N184_O) );
buf1 gate1236( .a(N185_I), .O(N185_O) );
buf1 gate1237( .a(N186_I), .O(N186_O) );
buf1 gate1238( .a(N187_I), .O(N187_O) );
buf1 gate1239( .a(N188_I), .O(N188_O) );
buf1 gate1240( .a(N189_I), .O(N189_O) );
buf1 gate1241( .a(N190_I), .O(N190_O) );
buf1 gate1242( .a(N191_I), .O(N191_O) );
buf1 gate1243( .a(N192_I), .O(N192_O) );
buf1 gate1244( .a(N193_I), .O(N193_O) );
buf1 gate1245( .a(N194_I), .O(N194_O) );
buf1 gate1246( .a(N195_I), .O(N195_O) );
buf1 gate1247( .a(N196_I), .O(N196_O) );
buf1 gate1248( .a(N197_I), .O(N197_O) );
buf1 gate1249( .a(N198_I), .O(N198_O) );
buf1 gate1250( .a(N199_I), .O(N199_O) );
buf1 gate1251( .a(N200_I), .O(N200_O) );
buf1 gate1252( .a(N201_I), .O(N201_O) );
buf1 gate1253( .a(N202_I), .O(N202_O) );
buf1 gate1254( .a(N203_I), .O(N203_O) );
buf1 gate1255( .a(N204_I), .O(N204_O) );
buf1 gate1256( .a(N205_I), .O(N205_O) );
buf1 gate1257( .a(N206_I), .O(N206_O) );
buf1 gate1258( .a(N207_I), .O(N207_O) );
buf1 gate1259( .a(N208_I), .O(N208_O) );
buf1 gate1260( .a(N209_I), .O(N209_O) );
buf1 gate1261( .a(N210_I), .O(N210_O) );
buf1 gate1262( .a(N211_I), .O(N211_O) );
buf1 gate1263( .a(N212_I), .O(N212_O) );
buf1 gate1264( .a(N213_I), .O(N213_O) );
buf1 gate1265( .a(N214_I), .O(N214_O) );
buf1 gate1266( .a(N215_I), .O(N215_O) );
buf1 gate1267( .a(N216_I), .O(N216_O) );
buf1 gate1268( .a(N217_I), .O(N217_O) );
buf1 gate1269( .a(N218_I), .O(N218_O) );

endmodule